module router 
(
  clk, 
  creditin_0, 
  creditin_1, 
  currx, 
  curry, 
  flitin_0, 
  flitin_1, 
  reset, 
  seu, 
  creditout_0,
  creditout_1,
  flitout_0,
  flitout_1
);
  input clk;
  input creditin_0;
  input creditin_1;
  input [2:0] currx;
  input [2:0] curry;
  input [11:0] flitin_0;
  input [11:0] flitin_1;
  input reset;
  input seu;
  output creditout_0;
  output creditout_1;
  output [11:0] flitout_0;
  output [11:0] flitout_1;
  wire c0nm__logic0_;
  wire c0nm_b0m__logic0_;
  wire c0nm_b0m_dqenablereg;
  wire c0nm_b0m_headflit_10_;
  wire c0nm_b0m_headflit_11_;
  wire c0nm_b0m_headflit_8_;
  wire c0nm_b0m_headflit_9_;
  wire c0nm_b0m_n1;
  wire c0nm_b0m_n9;
  wire [11:0] c0nm_b0m_rdata;
  wire c0nm_b0m_v0m_buffers0_0_;
  wire c0nm_b0m_v0m_buffers0_10_;
  wire c0nm_b0m_v0m_buffers0_11_;
  wire c0nm_b0m_v0m_buffers0_1_;
  wire c0nm_b0m_v0m_buffers0_2_;
  wire c0nm_b0m_v0m_buffers0_3_;
  wire c0nm_b0m_v0m_buffers0_4_;
  wire c0nm_b0m_v0m_buffers0_5_;
  wire c0nm_b0m_v0m_buffers0_6_;
  wire c0nm_b0m_v0m_buffers0_7_;
  wire c0nm_b0m_v0m_buffers0_8_;
  wire c0nm_b0m_v0m_buffers0_9_;
  wire c0nm_b0m_v0m_buffers2_0_;
  wire c0nm_b0m_v0m_buffers2_10_;
  wire c0nm_b0m_v0m_buffers2_11_;
  wire c0nm_b0m_v0m_buffers2_1_;
  wire c0nm_b0m_v0m_buffers2_2_;
  wire c0nm_b0m_v0m_buffers2_3_;
  wire c0nm_b0m_v0m_buffers2_4_;
  wire c0nm_b0m_v0m_buffers2_5_;
  wire c0nm_b0m_v0m_buffers2_6_;
  wire c0nm_b0m_v0m_buffers2_7_;
  wire c0nm_b0m_v0m_buffers2_8_;
  wire c0nm_b0m_v0m_buffers2_9_;
  wire c0nm_b0m_v0m_buffers3_0_;
  wire c0nm_b0m_v0m_buffers3_10_;
  wire c0nm_b0m_v0m_buffers3_11_;
  wire c0nm_b0m_v0m_buffers3_1_;
  wire c0nm_b0m_v0m_buffers3_2_;
  wire c0nm_b0m_v0m_buffers3_3_;
  wire c0nm_b0m_v0m_buffers3_4_;
  wire c0nm_b0m_v0m_buffers3_5_;
  wire c0nm_b0m_v0m_buffers3_6_;
  wire c0nm_b0m_v0m_buffers3_7_;
  wire c0nm_b0m_v0m_buffers3_8_;
  wire c0nm_b0m_v0m_buffers3_9_;
  wire c0nm_b0m_v0m_head_0_;
  wire c0nm_b0m_v0m_head_1_;
  wire c0nm_b0m_v0m_head_2_;
  wire c0nm_b0m_v0m_n1;
  wire c0nm_b0m_v0m_n10;
  wire c0nm_b0m_v0m_n100;
  wire c0nm_b0m_v0m_n101;
  wire c0nm_b0m_v0m_n102;
  wire c0nm_b0m_v0m_n103;
  wire c0nm_b0m_v0m_n104;
  wire c0nm_b0m_v0m_n105;
  wire c0nm_b0m_v0m_n106;
  wire c0nm_b0m_v0m_n107;
  wire c0nm_b0m_v0m_n108;
  wire c0nm_b0m_v0m_n109;
  wire c0nm_b0m_v0m_n11;
  wire c0nm_b0m_v0m_n110;
  wire c0nm_b0m_v0m_n111;
  wire c0nm_b0m_v0m_n112;
  wire c0nm_b0m_v0m_n113;
  wire c0nm_b0m_v0m_n114;
  wire c0nm_b0m_v0m_n115;
  wire c0nm_b0m_v0m_n116;
  wire c0nm_b0m_v0m_n117;
  wire c0nm_b0m_v0m_n118;
  wire c0nm_b0m_v0m_n119;
  wire c0nm_b0m_v0m_n12;
  wire c0nm_b0m_v0m_n120;
  wire c0nm_b0m_v0m_n121;
  wire c0nm_b0m_v0m_n122;
  wire c0nm_b0m_v0m_n123;
  wire c0nm_b0m_v0m_n124;
  wire c0nm_b0m_v0m_n125;
  wire c0nm_b0m_v0m_n126;
  wire c0nm_b0m_v0m_n127;
  wire c0nm_b0m_v0m_n128;
  wire c0nm_b0m_v0m_n129;
  wire c0nm_b0m_v0m_n13;
  wire c0nm_b0m_v0m_n130;
  wire c0nm_b0m_v0m_n131;
  wire c0nm_b0m_v0m_n132;
  wire c0nm_b0m_v0m_n133;
  wire c0nm_b0m_v0m_n134;
  wire c0nm_b0m_v0m_n135;
  wire c0nm_b0m_v0m_n136;
  wire c0nm_b0m_v0m_n137;
  wire c0nm_b0m_v0m_n138;
  wire c0nm_b0m_v0m_n139;
  wire c0nm_b0m_v0m_n14;
  wire c0nm_b0m_v0m_n140;
  wire c0nm_b0m_v0m_n141;
  wire c0nm_b0m_v0m_n142;
  wire c0nm_b0m_v0m_n143;
  wire c0nm_b0m_v0m_n144;
  wire c0nm_b0m_v0m_n145;
  wire c0nm_b0m_v0m_n146;
  wire c0nm_b0m_v0m_n147;
  wire c0nm_b0m_v0m_n148;
  wire c0nm_b0m_v0m_n149;
  wire c0nm_b0m_v0m_n15;
  wire c0nm_b0m_v0m_n150;
  wire c0nm_b0m_v0m_n151;
  wire c0nm_b0m_v0m_n152;
  wire c0nm_b0m_v0m_n153;
  wire c0nm_b0m_v0m_n154;
  wire c0nm_b0m_v0m_n155;
  wire c0nm_b0m_v0m_n156;
  wire c0nm_b0m_v0m_n157;
  wire c0nm_b0m_v0m_n158;
  wire c0nm_b0m_v0m_n159;
  wire c0nm_b0m_v0m_n16;
  wire c0nm_b0m_v0m_n160;
  wire c0nm_b0m_v0m_n161;
  wire c0nm_b0m_v0m_n162;
  wire c0nm_b0m_v0m_n163;
  wire c0nm_b0m_v0m_n164;
  wire c0nm_b0m_v0m_n165;
  wire c0nm_b0m_v0m_n166;
  wire c0nm_b0m_v0m_n167;
  wire c0nm_b0m_v0m_n168;
  wire c0nm_b0m_v0m_n169;
  wire c0nm_b0m_v0m_n17;
  wire c0nm_b0m_v0m_n170;
  wire c0nm_b0m_v0m_n171;
  wire c0nm_b0m_v0m_n1710;
  wire c0nm_b0m_v0m_n172;
  wire c0nm_b0m_v0m_n173;
  wire c0nm_b0m_v0m_n174;
  wire c0nm_b0m_v0m_n175;
  wire c0nm_b0m_v0m_n176;
  wire c0nm_b0m_v0m_n177;
  wire c0nm_b0m_v0m_n178;
  wire c0nm_b0m_v0m_n179;
  wire c0nm_b0m_v0m_n18;
  wire c0nm_b0m_v0m_n180;
  wire c0nm_b0m_v0m_n181;
  wire c0nm_b0m_v0m_n182;
  wire c0nm_b0m_v0m_n183;
  wire c0nm_b0m_v0m_n184;
  wire c0nm_b0m_v0m_n185;
  wire c0nm_b0m_v0m_n186;
  wire c0nm_b0m_v0m_n187;
  wire c0nm_b0m_v0m_n188;
  wire c0nm_b0m_v0m_n189;
  wire c0nm_b0m_v0m_n19;
  wire c0nm_b0m_v0m_n190;
  wire c0nm_b0m_v0m_n192;
  wire c0nm_b0m_v0m_n193;
  wire c0nm_b0m_v0m_n194;
  wire c0nm_b0m_v0m_n195;
  wire c0nm_b0m_v0m_n196;
  wire c0nm_b0m_v0m_n197;
  wire c0nm_b0m_v0m_n198;
  wire c0nm_b0m_v0m_n199;
  wire c0nm_b0m_v0m_n2;
  wire c0nm_b0m_v0m_n20;
  wire c0nm_b0m_v0m_n200;
  wire c0nm_b0m_v0m_n201;
  wire c0nm_b0m_v0m_n202;
  wire c0nm_b0m_v0m_n203;
  wire c0nm_b0m_v0m_n204;
  wire c0nm_b0m_v0m_n205;
  wire c0nm_b0m_v0m_n206;
  wire c0nm_b0m_v0m_n207;
  wire c0nm_b0m_v0m_n208;
  wire c0nm_b0m_v0m_n209;
  wire c0nm_b0m_v0m_n21;
  wire c0nm_b0m_v0m_n210;
  wire c0nm_b0m_v0m_n211;
  wire c0nm_b0m_v0m_n212;
  wire c0nm_b0m_v0m_n213;
  wire c0nm_b0m_v0m_n214;
  wire c0nm_b0m_v0m_n215;
  wire c0nm_b0m_v0m_n216;
  wire c0nm_b0m_v0m_n217;
  wire c0nm_b0m_v0m_n218;
  wire c0nm_b0m_v0m_n219;
  wire c0nm_b0m_v0m_n22;
  wire c0nm_b0m_v0m_n220;
  wire c0nm_b0m_v0m_n221;
  wire c0nm_b0m_v0m_n222;
  wire c0nm_b0m_v0m_n223;
  wire c0nm_b0m_v0m_n224;
  wire c0nm_b0m_v0m_n225;
  wire c0nm_b0m_v0m_n226;
  wire c0nm_b0m_v0m_n227;
  wire c0nm_b0m_v0m_n228;
  wire c0nm_b0m_v0m_n229;
  wire c0nm_b0m_v0m_n23;
  wire c0nm_b0m_v0m_n230;
  wire c0nm_b0m_v0m_n231;
  wire c0nm_b0m_v0m_n232;
  wire c0nm_b0m_v0m_n233;
  wire c0nm_b0m_v0m_n234;
  wire c0nm_b0m_v0m_n235;
  wire c0nm_b0m_v0m_n236;
  wire c0nm_b0m_v0m_n237;
  wire c0nm_b0m_v0m_n238;
  wire c0nm_b0m_v0m_n239;
  wire c0nm_b0m_v0m_n24;
  wire c0nm_b0m_v0m_n240;
  wire c0nm_b0m_v0m_n241;
  wire c0nm_b0m_v0m_n242;
  wire c0nm_b0m_v0m_n243;
  wire c0nm_b0m_v0m_n244;
  wire c0nm_b0m_v0m_n245;
  wire c0nm_b0m_v0m_n246;
  wire c0nm_b0m_v0m_n247;
  wire c0nm_b0m_v0m_n248;
  wire c0nm_b0m_v0m_n249;
  wire c0nm_b0m_v0m_n25;
  wire c0nm_b0m_v0m_n250;
  wire c0nm_b0m_v0m_n251;
  wire c0nm_b0m_v0m_n252;
  wire c0nm_b0m_v0m_n253;
  wire c0nm_b0m_v0m_n254;
  wire c0nm_b0m_v0m_n255;
  wire c0nm_b0m_v0m_n256;
  wire c0nm_b0m_v0m_n257;
  wire c0nm_b0m_v0m_n258;
  wire c0nm_b0m_v0m_n259;
  wire c0nm_b0m_v0m_n26;
  wire c0nm_b0m_v0m_n260;
  wire c0nm_b0m_v0m_n261;
  wire c0nm_b0m_v0m_n262;
  wire c0nm_b0m_v0m_n263;
  wire c0nm_b0m_v0m_n264;
  wire c0nm_b0m_v0m_n265;
  wire c0nm_b0m_v0m_n266;
  wire c0nm_b0m_v0m_n267;
  wire c0nm_b0m_v0m_n268;
  wire c0nm_b0m_v0m_n269;
  wire c0nm_b0m_v0m_n27;
  wire c0nm_b0m_v0m_n270;
  wire c0nm_b0m_v0m_n271;
  wire c0nm_b0m_v0m_n272;
  wire c0nm_b0m_v0m_n273;
  wire c0nm_b0m_v0m_n274;
  wire c0nm_b0m_v0m_n275;
  wire c0nm_b0m_v0m_n276;
  wire c0nm_b0m_v0m_n28;
  wire c0nm_b0m_v0m_n29;
  wire c0nm_b0m_v0m_n3;
  wire c0nm_b0m_v0m_n30;
  wire c0nm_b0m_v0m_n31;
  wire c0nm_b0m_v0m_n32;
  wire c0nm_b0m_v0m_n33;
  wire c0nm_b0m_v0m_n34;
  wire c0nm_b0m_v0m_n35;
  wire c0nm_b0m_v0m_n36;
  wire c0nm_b0m_v0m_n37;
  wire c0nm_b0m_v0m_n38;
  wire c0nm_b0m_v0m_n39;
  wire c0nm_b0m_v0m_n4;
  wire c0nm_b0m_v0m_n40;
  wire c0nm_b0m_v0m_n41;
  wire c0nm_b0m_v0m_n42;
  wire c0nm_b0m_v0m_n43;
  wire c0nm_b0m_v0m_n44;
  wire c0nm_b0m_v0m_n45;
  wire c0nm_b0m_v0m_n46;
  wire c0nm_b0m_v0m_n47;
  wire c0nm_b0m_v0m_n48;
  wire c0nm_b0m_v0m_n49;
  wire c0nm_b0m_v0m_n5;
  wire c0nm_b0m_v0m_n50;
  wire c0nm_b0m_v0m_n51;
  wire c0nm_b0m_v0m_n52;
  wire c0nm_b0m_v0m_n53;
  wire c0nm_b0m_v0m_n54;
  wire c0nm_b0m_v0m_n55;
  wire c0nm_b0m_v0m_n56;
  wire c0nm_b0m_v0m_n57;
  wire c0nm_b0m_v0m_n58;
  wire c0nm_b0m_v0m_n59;
  wire c0nm_b0m_v0m_n6;
  wire c0nm_b0m_v0m_n60;
  wire c0nm_b0m_v0m_n61;
  wire c0nm_b0m_v0m_n62;
  wire c0nm_b0m_v0m_n63;
  wire c0nm_b0m_v0m_n64;
  wire c0nm_b0m_v0m_n65;
  wire c0nm_b0m_v0m_n66;
  wire c0nm_b0m_v0m_n67;
  wire c0nm_b0m_v0m_n68;
  wire c0nm_b0m_v0m_n69;
  wire c0nm_b0m_v0m_n7;
  wire c0nm_b0m_v0m_n70;
  wire c0nm_b0m_v0m_n71;
  wire c0nm_b0m_v0m_n72;
  wire c0nm_b0m_v0m_n73;
  wire c0nm_b0m_v0m_n74;
  wire c0nm_b0m_v0m_n75;
  wire c0nm_b0m_v0m_n76;
  wire c0nm_b0m_v0m_n77;
  wire c0nm_b0m_v0m_n78;
  wire c0nm_b0m_v0m_n79;
  wire c0nm_b0m_v0m_n8;
  wire c0nm_b0m_v0m_n80;
  wire c0nm_b0m_v0m_n81;
  wire c0nm_b0m_v0m_n82;
  wire c0nm_b0m_v0m_n83;
  wire c0nm_b0m_v0m_n84;
  wire c0nm_b0m_v0m_n85;
  wire c0nm_b0m_v0m_n86;
  wire c0nm_b0m_v0m_n87;
  wire c0nm_b0m_v0m_n88;
  wire c0nm_b0m_v0m_n89;
  wire c0nm_b0m_v0m_n9;
  wire c0nm_b0m_v0m_n90;
  wire c0nm_b0m_v0m_n91;
  wire c0nm_b0m_v0m_n92;
  wire c0nm_b0m_v0m_n93;
  wire c0nm_b0m_v0m_n94;
  wire c0nm_b0m_v0m_n95;
  wire c0nm_b0m_v0m_n96;
  wire c0nm_b0m_v0m_n97;
  wire c0nm_b0m_v0m_n98;
  wire c0nm_b0m_v0m_n99;
  wire c0nm_b0m_v0m_tail_0_;
  wire c0nm_b0m_v0m_tail_1_;
  wire c0nm_b0m_wdata_10_;
  wire c0nm_b0m_wdata_11_;
  wire c0nm_b0m_wdata_2_;
  wire c0nm_b0m_wdata_3_;
  wire c0nm_b0m_wdata_4_;
  wire c0nm_b0m_wdata_5_;
  wire c0nm_b0m_wdata_6_;
  wire c0nm_b0m_wdata_7_;
  wire c0nm_b0m_wdata_8_;
  wire c0nm_b0m_wdata_9_;
  wire [7:0] c0nm_headflit;
  wire c0nm_n1;
  wire c0nm_n2;
  wire c0nm_r0m_n1;
  wire c0nm_r0m_n10;
  wire c0nm_r0m_n100;
  wire c0nm_r0m_n11;
  wire c0nm_r0m_n110;
  wire c0nm_r0m_n12;
  wire c0nm_r0m_n13;
  wire c0nm_r0m_n14;
  wire c0nm_r0m_n15;
  wire c0nm_r0m_n16;
  wire c0nm_r0m_n2;
  wire c0nm_r0m_n3;
  wire c0nm_r0m_n4;
  wire c0nm_r0m_n5;
  wire c0nm_r0m_n6;
  wire c0nm_r0m_n7;
  wire c0nm_r0m_n8;
  wire c0nm_r0m_n9;
  wire [1:0] c0nm_routewire;
  wire c0nm_v0m_full;
  wire c0nm_v0m_n1;
  wire c0nm_v0m_n10;
  wire c0nm_v0m_n11;
  wire c0nm_v0m_n12;
  wire c0nm_v0m_n13;
  wire c0nm_v0m_n14;
  wire c0nm_v0m_n15;
  wire c0nm_v0m_n16;
  wire c0nm_v0m_n17;
  wire c0nm_v0m_n18;
  wire c0nm_v0m_n19;
  wire c0nm_v0m_n2;
  wire c0nm_v0m_n20;
  wire c0nm_v0m_n21;
  wire c0nm_v0m_n22;
  wire c0nm_v0m_n23;
  wire c0nm_v0m_n24;
  wire c0nm_v0m_n25;
  wire c0nm_v0m_n26;
  wire c0nm_v0m_n27;
  wire c0nm_v0m_n28;
  wire c0nm_v0m_n29;
  wire c0nm_v0m_n3;
  wire c0nm_v0m_n30;
  wire c0nm_v0m_n31;
  wire c0nm_v0m_n4;
  wire c0nm_v0m_n5;
  wire c0nm_v0m_n57;
  wire c0nm_v0m_n58;
  wire c0nm_v0m_n6;
  wire c0nm_v0m_n61;
  wire c0nm_v0m_n62;
  wire c0nm_v0m_n63;
  wire c0nm_v0m_n64;
  wire c0nm_v0m_n7;
  wire c0nm_v0m_n8;
  wire c0nm_v0m_n9;
  wire c0nm_v0m_state_queuelen_0_;
  wire c0nm_v0m_state_queuelen_1_;
  wire c0nm_v0m_state_queuelen_2_;
  wire c0nm_v0m_state_status_0_;
  wire c0nm_v0m_state_status_1_;
  wire c0sm__logic0_;
  wire c0sm_b0m__logic0_;
  wire c0sm_b0m_dqenablereg;
  wire c0sm_b0m_headflit_10_;
  wire c0sm_b0m_headflit_11_;
  wire c0sm_b0m_headflit_8_;
  wire c0sm_b0m_headflit_9_;
  wire c0sm_b0m_n2;
  wire c0sm_b0m_n9;
  wire [11:0] c0sm_b0m_rdata;
  wire c0sm_b0m_v0m_buffers0_0_;
  wire c0sm_b0m_v0m_buffers0_10_;
  wire c0sm_b0m_v0m_buffers0_11_;
  wire c0sm_b0m_v0m_buffers0_1_;
  wire c0sm_b0m_v0m_buffers0_2_;
  wire c0sm_b0m_v0m_buffers0_3_;
  wire c0sm_b0m_v0m_buffers0_4_;
  wire c0sm_b0m_v0m_buffers0_5_;
  wire c0sm_b0m_v0m_buffers0_6_;
  wire c0sm_b0m_v0m_buffers0_7_;
  wire c0sm_b0m_v0m_buffers0_8_;
  wire c0sm_b0m_v0m_buffers0_9_;
  wire c0sm_b0m_v0m_buffers2_0_;
  wire c0sm_b0m_v0m_buffers2_10_;
  wire c0sm_b0m_v0m_buffers2_11_;
  wire c0sm_b0m_v0m_buffers2_1_;
  wire c0sm_b0m_v0m_buffers2_2_;
  wire c0sm_b0m_v0m_buffers2_3_;
  wire c0sm_b0m_v0m_buffers2_4_;
  wire c0sm_b0m_v0m_buffers2_5_;
  wire c0sm_b0m_v0m_buffers2_6_;
  wire c0sm_b0m_v0m_buffers2_7_;
  wire c0sm_b0m_v0m_buffers2_8_;
  wire c0sm_b0m_v0m_buffers2_9_;
  wire c0sm_b0m_v0m_buffers3_0_;
  wire c0sm_b0m_v0m_buffers3_10_;
  wire c0sm_b0m_v0m_buffers3_11_;
  wire c0sm_b0m_v0m_buffers3_1_;
  wire c0sm_b0m_v0m_buffers3_2_;
  wire c0sm_b0m_v0m_buffers3_3_;
  wire c0sm_b0m_v0m_buffers3_4_;
  wire c0sm_b0m_v0m_buffers3_5_;
  wire c0sm_b0m_v0m_buffers3_6_;
  wire c0sm_b0m_v0m_buffers3_7_;
  wire c0sm_b0m_v0m_buffers3_8_;
  wire c0sm_b0m_v0m_buffers3_9_;
  wire c0sm_b0m_v0m_head_0_;
  wire c0sm_b0m_v0m_head_1_;
  wire c0sm_b0m_v0m_head_2_;
  wire c0sm_b0m_v0m_n1;
  wire c0sm_b0m_v0m_n10;
  wire c0sm_b0m_v0m_n100;
  wire c0sm_b0m_v0m_n101;
  wire c0sm_b0m_v0m_n102;
  wire c0sm_b0m_v0m_n103;
  wire c0sm_b0m_v0m_n104;
  wire c0sm_b0m_v0m_n105;
  wire c0sm_b0m_v0m_n106;
  wire c0sm_b0m_v0m_n107;
  wire c0sm_b0m_v0m_n108;
  wire c0sm_b0m_v0m_n109;
  wire c0sm_b0m_v0m_n11;
  wire c0sm_b0m_v0m_n110;
  wire c0sm_b0m_v0m_n111;
  wire c0sm_b0m_v0m_n112;
  wire c0sm_b0m_v0m_n113;
  wire c0sm_b0m_v0m_n114;
  wire c0sm_b0m_v0m_n115;
  wire c0sm_b0m_v0m_n116;
  wire c0sm_b0m_v0m_n117;
  wire c0sm_b0m_v0m_n118;
  wire c0sm_b0m_v0m_n119;
  wire c0sm_b0m_v0m_n12;
  wire c0sm_b0m_v0m_n120;
  wire c0sm_b0m_v0m_n121;
  wire c0sm_b0m_v0m_n122;
  wire c0sm_b0m_v0m_n123;
  wire c0sm_b0m_v0m_n124;
  wire c0sm_b0m_v0m_n125;
  wire c0sm_b0m_v0m_n126;
  wire c0sm_b0m_v0m_n127;
  wire c0sm_b0m_v0m_n128;
  wire c0sm_b0m_v0m_n129;
  wire c0sm_b0m_v0m_n13;
  wire c0sm_b0m_v0m_n130;
  wire c0sm_b0m_v0m_n131;
  wire c0sm_b0m_v0m_n132;
  wire c0sm_b0m_v0m_n133;
  wire c0sm_b0m_v0m_n134;
  wire c0sm_b0m_v0m_n135;
  wire c0sm_b0m_v0m_n136;
  wire c0sm_b0m_v0m_n137;
  wire c0sm_b0m_v0m_n138;
  wire c0sm_b0m_v0m_n139;
  wire c0sm_b0m_v0m_n14;
  wire c0sm_b0m_v0m_n140;
  wire c0sm_b0m_v0m_n141;
  wire c0sm_b0m_v0m_n142;
  wire c0sm_b0m_v0m_n143;
  wire c0sm_b0m_v0m_n144;
  wire c0sm_b0m_v0m_n145;
  wire c0sm_b0m_v0m_n146;
  wire c0sm_b0m_v0m_n147;
  wire c0sm_b0m_v0m_n148;
  wire c0sm_b0m_v0m_n149;
  wire c0sm_b0m_v0m_n15;
  wire c0sm_b0m_v0m_n150;
  wire c0sm_b0m_v0m_n151;
  wire c0sm_b0m_v0m_n152;
  wire c0sm_b0m_v0m_n153;
  wire c0sm_b0m_v0m_n154;
  wire c0sm_b0m_v0m_n155;
  wire c0sm_b0m_v0m_n156;
  wire c0sm_b0m_v0m_n157;
  wire c0sm_b0m_v0m_n158;
  wire c0sm_b0m_v0m_n159;
  wire c0sm_b0m_v0m_n16;
  wire c0sm_b0m_v0m_n160;
  wire c0sm_b0m_v0m_n161;
  wire c0sm_b0m_v0m_n162;
  wire c0sm_b0m_v0m_n163;
  wire c0sm_b0m_v0m_n164;
  wire c0sm_b0m_v0m_n165;
  wire c0sm_b0m_v0m_n166;
  wire c0sm_b0m_v0m_n167;
  wire c0sm_b0m_v0m_n168;
  wire c0sm_b0m_v0m_n169;
  wire c0sm_b0m_v0m_n17;
  wire c0sm_b0m_v0m_n170;
  wire c0sm_b0m_v0m_n171;
  wire c0sm_b0m_v0m_n1710;
  wire c0sm_b0m_v0m_n172;
  wire c0sm_b0m_v0m_n173;
  wire c0sm_b0m_v0m_n174;
  wire c0sm_b0m_v0m_n175;
  wire c0sm_b0m_v0m_n176;
  wire c0sm_b0m_v0m_n177;
  wire c0sm_b0m_v0m_n178;
  wire c0sm_b0m_v0m_n179;
  wire c0sm_b0m_v0m_n18;
  wire c0sm_b0m_v0m_n180;
  wire c0sm_b0m_v0m_n181;
  wire c0sm_b0m_v0m_n182;
  wire c0sm_b0m_v0m_n183;
  wire c0sm_b0m_v0m_n184;
  wire c0sm_b0m_v0m_n185;
  wire c0sm_b0m_v0m_n186;
  wire c0sm_b0m_v0m_n187;
  wire c0sm_b0m_v0m_n188;
  wire c0sm_b0m_v0m_n189;
  wire c0sm_b0m_v0m_n19;
  wire c0sm_b0m_v0m_n190;
  wire c0sm_b0m_v0m_n192;
  wire c0sm_b0m_v0m_n193;
  wire c0sm_b0m_v0m_n194;
  wire c0sm_b0m_v0m_n195;
  wire c0sm_b0m_v0m_n2;
  wire c0sm_b0m_v0m_n20;
  wire c0sm_b0m_v0m_n21;
  wire c0sm_b0m_v0m_n22;
  wire c0sm_b0m_v0m_n23;
  wire c0sm_b0m_v0m_n24;
  wire c0sm_b0m_v0m_n25;
  wire c0sm_b0m_v0m_n26;
  wire c0sm_b0m_v0m_n262;
  wire c0sm_b0m_v0m_n263;
  wire c0sm_b0m_v0m_n264;
  wire c0sm_b0m_v0m_n265;
  wire c0sm_b0m_v0m_n266;
  wire c0sm_b0m_v0m_n267;
  wire c0sm_b0m_v0m_n268;
  wire c0sm_b0m_v0m_n269;
  wire c0sm_b0m_v0m_n27;
  wire c0sm_b0m_v0m_n270;
  wire c0sm_b0m_v0m_n271;
  wire c0sm_b0m_v0m_n272;
  wire c0sm_b0m_v0m_n273;
  wire c0sm_b0m_v0m_n274;
  wire c0sm_b0m_v0m_n275;
  wire c0sm_b0m_v0m_n276;
  wire c0sm_b0m_v0m_n277;
  wire c0sm_b0m_v0m_n278;
  wire c0sm_b0m_v0m_n279;
  wire c0sm_b0m_v0m_n28;
  wire c0sm_b0m_v0m_n280;
  wire c0sm_b0m_v0m_n281;
  wire c0sm_b0m_v0m_n282;
  wire c0sm_b0m_v0m_n283;
  wire c0sm_b0m_v0m_n284;
  wire c0sm_b0m_v0m_n285;
  wire c0sm_b0m_v0m_n286;
  wire c0sm_b0m_v0m_n287;
  wire c0sm_b0m_v0m_n288;
  wire c0sm_b0m_v0m_n289;
  wire c0sm_b0m_v0m_n29;
  wire c0sm_b0m_v0m_n290;
  wire c0sm_b0m_v0m_n291;
  wire c0sm_b0m_v0m_n292;
  wire c0sm_b0m_v0m_n293;
  wire c0sm_b0m_v0m_n294;
  wire c0sm_b0m_v0m_n295;
  wire c0sm_b0m_v0m_n296;
  wire c0sm_b0m_v0m_n297;
  wire c0sm_b0m_v0m_n298;
  wire c0sm_b0m_v0m_n299;
  wire c0sm_b0m_v0m_n3;
  wire c0sm_b0m_v0m_n30;
  wire c0sm_b0m_v0m_n300;
  wire c0sm_b0m_v0m_n301;
  wire c0sm_b0m_v0m_n302;
  wire c0sm_b0m_v0m_n303;
  wire c0sm_b0m_v0m_n304;
  wire c0sm_b0m_v0m_n305;
  wire c0sm_b0m_v0m_n306;
  wire c0sm_b0m_v0m_n307;
  wire c0sm_b0m_v0m_n308;
  wire c0sm_b0m_v0m_n309;
  wire c0sm_b0m_v0m_n31;
  wire c0sm_b0m_v0m_n310;
  wire c0sm_b0m_v0m_n311;
  wire c0sm_b0m_v0m_n312;
  wire c0sm_b0m_v0m_n313;
  wire c0sm_b0m_v0m_n314;
  wire c0sm_b0m_v0m_n315;
  wire c0sm_b0m_v0m_n316;
  wire c0sm_b0m_v0m_n317;
  wire c0sm_b0m_v0m_n318;
  wire c0sm_b0m_v0m_n319;
  wire c0sm_b0m_v0m_n32;
  wire c0sm_b0m_v0m_n320;
  wire c0sm_b0m_v0m_n321;
  wire c0sm_b0m_v0m_n322;
  wire c0sm_b0m_v0m_n323;
  wire c0sm_b0m_v0m_n324;
  wire c0sm_b0m_v0m_n325;
  wire c0sm_b0m_v0m_n326;
  wire c0sm_b0m_v0m_n327;
  wire c0sm_b0m_v0m_n328;
  wire c0sm_b0m_v0m_n329;
  wire c0sm_b0m_v0m_n33;
  wire c0sm_b0m_v0m_n330;
  wire c0sm_b0m_v0m_n331;
  wire c0sm_b0m_v0m_n332;
  wire c0sm_b0m_v0m_n333;
  wire c0sm_b0m_v0m_n334;
  wire c0sm_b0m_v0m_n335;
  wire c0sm_b0m_v0m_n336;
  wire c0sm_b0m_v0m_n337;
  wire c0sm_b0m_v0m_n338;
  wire c0sm_b0m_v0m_n339;
  wire c0sm_b0m_v0m_n34;
  wire c0sm_b0m_v0m_n340;
  wire c0sm_b0m_v0m_n341;
  wire c0sm_b0m_v0m_n342;
  wire c0sm_b0m_v0m_n343;
  wire c0sm_b0m_v0m_n344;
  wire c0sm_b0m_v0m_n345;
  wire c0sm_b0m_v0m_n346;
  wire c0sm_b0m_v0m_n347;
  wire c0sm_b0m_v0m_n348;
  wire c0sm_b0m_v0m_n349;
  wire c0sm_b0m_v0m_n35;
  wire c0sm_b0m_v0m_n350;
  wire c0sm_b0m_v0m_n351;
  wire c0sm_b0m_v0m_n352;
  wire c0sm_b0m_v0m_n353;
  wire c0sm_b0m_v0m_n354;
  wire c0sm_b0m_v0m_n355;
  wire c0sm_b0m_v0m_n36;
  wire c0sm_b0m_v0m_n37;
  wire c0sm_b0m_v0m_n38;
  wire c0sm_b0m_v0m_n39;
  wire c0sm_b0m_v0m_n40;
  wire c0sm_b0m_v0m_n41;
  wire c0sm_b0m_v0m_n42;
  wire c0sm_b0m_v0m_n43;
  wire c0sm_b0m_v0m_n44;
  wire c0sm_b0m_v0m_n45;
  wire c0sm_b0m_v0m_n46;
  wire c0sm_b0m_v0m_n47;
  wire c0sm_b0m_v0m_n48;
  wire c0sm_b0m_v0m_n49;
  wire c0sm_b0m_v0m_n5;
  wire c0sm_b0m_v0m_n6;
  wire c0sm_b0m_v0m_n62;
  wire c0sm_b0m_v0m_n63;
  wire c0sm_b0m_v0m_n64;
  wire c0sm_b0m_v0m_n65;
  wire c0sm_b0m_v0m_n66;
  wire c0sm_b0m_v0m_n67;
  wire c0sm_b0m_v0m_n68;
  wire c0sm_b0m_v0m_n69;
  wire c0sm_b0m_v0m_n7;
  wire c0sm_b0m_v0m_n70;
  wire c0sm_b0m_v0m_n71;
  wire c0sm_b0m_v0m_n72;
  wire c0sm_b0m_v0m_n73;
  wire c0sm_b0m_v0m_n74;
  wire c0sm_b0m_v0m_n75;
  wire c0sm_b0m_v0m_n76;
  wire c0sm_b0m_v0m_n77;
  wire c0sm_b0m_v0m_n78;
  wire c0sm_b0m_v0m_n79;
  wire c0sm_b0m_v0m_n8;
  wire c0sm_b0m_v0m_n80;
  wire c0sm_b0m_v0m_n81;
  wire c0sm_b0m_v0m_n82;
  wire c0sm_b0m_v0m_n83;
  wire c0sm_b0m_v0m_n84;
  wire c0sm_b0m_v0m_n85;
  wire c0sm_b0m_v0m_n86;
  wire c0sm_b0m_v0m_n87;
  wire c0sm_b0m_v0m_n88;
  wire c0sm_b0m_v0m_n89;
  wire c0sm_b0m_v0m_n90;
  wire c0sm_b0m_v0m_n91;
  wire c0sm_b0m_v0m_n92;
  wire c0sm_b0m_v0m_n93;
  wire c0sm_b0m_v0m_n94;
  wire c0sm_b0m_v0m_n95;
  wire c0sm_b0m_v0m_n96;
  wire c0sm_b0m_v0m_n97;
  wire c0sm_b0m_v0m_n98;
  wire c0sm_b0m_v0m_n99;
  wire c0sm_b0m_v0m_tail_0_;
  wire c0sm_b0m_v0m_tail_1_;
  wire c0sm_b0m_wdata_10_;
  wire c0sm_b0m_wdata_11_;
  wire c0sm_b0m_wdata_2_;
  wire c0sm_b0m_wdata_3_;
  wire c0sm_b0m_wdata_4_;
  wire c0sm_b0m_wdata_5_;
  wire c0sm_b0m_wdata_6_;
  wire c0sm_b0m_wdata_7_;
  wire c0sm_b0m_wdata_8_;
  wire c0sm_b0m_wdata_9_;
  wire [7:0] c0sm_headflit;
  wire c0sm_n3;
  wire c0sm_n4;
  wire c0sm_r0m_n1;
  wire c0sm_r0m_n10;
  wire c0sm_r0m_n100;
  wire c0sm_r0m_n11;
  wire c0sm_r0m_n110;
  wire c0sm_r0m_n12;
  wire c0sm_r0m_n13;
  wire c0sm_r0m_n14;
  wire c0sm_r0m_n15;
  wire c0sm_r0m_n16;
  wire c0sm_r0m_n2;
  wire c0sm_r0m_n3;
  wire c0sm_r0m_n5;
  wire c0sm_r0m_n6;
  wire c0sm_r0m_n7;
  wire c0sm_r0m_n8;
  wire c0sm_r0m_n9;
  wire [1:0] c0sm_routewire;
  wire c0sm_v0m_full;
  wire c0sm_v0m_n1;
  wire c0sm_v0m_n10;
  wire c0sm_v0m_n11;
  wire c0sm_v0m_n12;
  wire c0sm_v0m_n13;
  wire c0sm_v0m_n14;
  wire c0sm_v0m_n15;
  wire c0sm_v0m_n16;
  wire c0sm_v0m_n17;
  wire c0sm_v0m_n18;
  wire c0sm_v0m_n19;
  wire c0sm_v0m_n2;
  wire c0sm_v0m_n20;
  wire c0sm_v0m_n21;
  wire c0sm_v0m_n22;
  wire c0sm_v0m_n23;
  wire c0sm_v0m_n24;
  wire c0sm_v0m_n25;
  wire c0sm_v0m_n26;
  wire c0sm_v0m_n27;
  wire c0sm_v0m_n28;
  wire c0sm_v0m_n29;
  wire c0sm_v0m_n3;
  wire c0sm_v0m_n32;
  wire c0sm_v0m_n33;
  wire c0sm_v0m_n4;
  wire c0sm_v0m_n5;
  wire c0sm_v0m_n57;
  wire c0sm_v0m_n58;
  wire c0sm_v0m_n6;
  wire c0sm_v0m_n61;
  wire c0sm_v0m_n62;
  wire c0sm_v0m_n63;
  wire c0sm_v0m_n64;
  wire c0sm_v0m_n7;
  wire c0sm_v0m_n8;
  wire c0sm_v0m_n9;
  wire c0sm_v0m_state_queuelen_0_;
  wire c0sm_v0m_state_queuelen_1_;
  wire c0sm_v0m_state_queuelen_2_;
  wire c0sm_v0m_state_status_0_;
  wire c0sm_v0m_state_status_1_;
  wire [1:0] colsel0;
  wire [1:0] colsel1;
  wire debitout_0;
  wire debitout_1;
  wire [11:0] flitout_switch_0;
  wire [11:0] flitout_switch_1;
  wire net1;
  wire nomorebufs_0;
  wire nomorebufs_1;
  wire s0m__logic0_;
  wire s0m_debit_outvc0;
  wire s0m_debit_outvc1;
  wire s0m_elig_0_;
  wire s0m_elig_1_;
  wire s0m_m0m_n1;
  wire s0m_m0m_n10;
  wire s0m_m0m_n2;
  wire s0m_m0m_n3;
  wire s0m_m0m_row1_0_;
  wire s0m_m1m_n1;
  wire s0m_m1m_n10;
  wire s0m_m1m_n2;
  wire s0m_m1m_n3;
  wire s0m_m1m_row1_0_;
  wire s0m_n1;
  wire s0m_n10;
  wire s0m_n11;
  wire s0m_n12;
  wire s0m_n13;
  wire s0m_n14;
  wire s0m_n15;
  wire s0m_n16;
  wire s0m_n17;
  wire s0m_n18;
  wire s0m_n19;
  wire s0m_n2;
  wire s0m_n20;
  wire s0m_n22;
  wire s0m_n23;
  wire s0m_n24;
  wire s0m_n25;
  wire s0m_n26;
  wire s0m_n3;
  wire s0m_n4;
  wire s0m_n5;
  wire s0m_n6;
  wire s0m_n7;
  wire s0m_n8;
  wire s0m_n9;
  wire s0m_no_bufs0;
  wire s0m_no_bufs1;
  wire s0m_o0nm_n1;
  wire s0m_o0nm_n11;
  wire s0m_o0nm_n12;
  wire s0m_o0nm_n13;
  wire s0m_o0nm_n14;
  wire s0m_o0nm_n15;
  wire s0m_o0nm_n16;
  wire s0m_o0nm_n17;
  wire s0m_o0nm_n18;
  wire s0m_o0nm_n19;
  wire s0m_o0nm_n2;
  wire s0m_o0nm_n20;
  wire s0m_o0nm_n21;
  wire s0m_o0nm_n22;
  wire s0m_o0nm_n23;
  wire s0m_o0nm_n24;
  wire s0m_o0nm_n25;
  wire s0m_o0nm_n3;
  wire s0m_o0nm_n30;
  wire s0m_o0nm_n31;
  wire s0m_o0nm_n35;
  wire s0m_o0nm_n36;
  wire s0m_o0nm_n37;
  wire s0m_o0nm_n38;
  wire s0m_o0nm_n4;
  wire s0m_o0nm_n41;
  wire s0m_o0nm_n42;
  wire s0m_o0nm_n5;
  wire s0m_o0nm_n6;
  wire s0m_o0nm_n7;
  wire s0m_o0nm_n9;
  wire s0m_o0nm_state_assigned;
  wire s0m_o0nm_state_credits_0_;
  wire s0m_o0nm_state_credits_1_;
  wire s0m_o0nm_state_credits_2_;
  wire s0m_o0sm_n1;
  wire s0m_o0sm_n11;
  wire s0m_o0sm_n12;
  wire s0m_o0sm_n13;
  wire s0m_o0sm_n14;
  wire s0m_o0sm_n15;
  wire s0m_o0sm_n16;
  wire s0m_o0sm_n17;
  wire s0m_o0sm_n18;
  wire s0m_o0sm_n19;
  wire s0m_o0sm_n2;
  wire s0m_o0sm_n20;
  wire s0m_o0sm_n21;
  wire s0m_o0sm_n22;
  wire s0m_o0sm_n23;
  wire s0m_o0sm_n24;
  wire s0m_o0sm_n25;
  wire s0m_o0sm_n26;
  wire s0m_o0sm_n27;
  wire s0m_o0sm_n3;
  wire s0m_o0sm_n35;
  wire s0m_o0sm_n36;
  wire s0m_o0sm_n37;
  wire s0m_o0sm_n38;
  wire s0m_o0sm_n4;
  wire s0m_o0sm_n41;
  wire s0m_o0sm_n42;
  wire s0m_o0sm_n5;
  wire s0m_o0sm_n6;
  wire s0m_o0sm_n7;
  wire s0m_o0sm_n9;
  wire s0m_o0sm_state_assigned;
  wire s0m_o0sm_state_credits_0_;
  wire s0m_o0sm_state_credits_1_;
  wire s0m_o0sm_state_credits_2_;
  wire s0m_outb0_0_;
  wire s0m_outb0_1_;
  wire s0m_outb1_0_;
  wire s0m_outb1_1_;
  wire [1:0] s0m_request0;
  wire [1:0] s0m_request1;
  wire s0m_state_invc0_0_;
  wire s0m_state_invc0_1_;
  wire s0m_state_invc1_0_;
  wire s0m_state_invc1_1_;
  wire s0m_tail_outvc0;
  wire s0m_tail_outvc1;
  wire [1:0] swalloc_req_0;
  wire [1:0] swalloc_req_1;
  wire [1:0] swalloc_resp_0;
  wire [1:0] swalloc_resp_1;
  wire tailout_0;
  wire tailout_1;
  wire x0m__logic0_;
  wire x0m__logic1_;
  wire x0m_bx0m_m0m_int01;
  wire x0m_bx0m_m1m_int01;
  wire x0m_bx10m_m0m_int01;
  wire x0m_bx10m_m1m_int01;
  wire x0m_bx11m_m0m_int01;
  wire x0m_bx11m_m1m_int01;
  wire x0m_bx1m_m0m_int01;
  wire x0m_bx1m_m1m_int01;
  wire x0m_bx2m_m0m_int01;
  wire x0m_bx2m_m1m_int01;
  wire x0m_bx3m_m0m_int01;
  wire x0m_bx3m_m1m_int01;
  wire x0m_bx4m_m0m_int01;
  wire x0m_bx4m_m1m_int01;
  wire x0m_bx5m_m0m_int01;
  wire x0m_bx5m_m1m_int01;
  wire x0m_bx6m_m0m_int01;
  wire x0m_bx6m_m1m_int01;
  wire x0m_bx7m_m0m_int01;
  wire x0m_bx7m_m1m_int01;
  wire x0m_bx8m_m0m_int01;
  wire x0m_bx8m_m1m_int01;
  wire x0m_bx9m_m0m_int01;
  wire x0m_bx9m_m1m_int01;
  wire x0m_colsel0reg_0_;
  wire x0m_colsel0reg_1_;
  wire x0m_colsel1reg_0_;
  wire x0m_colsel1reg_1_;
  wire x0m_n3;
  wire x0m_n4;
  wire x0m_n5;
  wire x0m_n6;
  // sz:2: index:0 c0nm_b0m_v0m_n262 c0nm_b0m_v0m_n263 
  // sz:2: index:1 c0nm_b0m_rdata[0] c0nm_b0m_rdata[1] 
  // sz:2: index:2 c0nm_b0m_v0m_n207 c0nm_b0m_v0m_n206 
  // sz:2: index:3 c0sm_b0m_v0m_n262 c0sm_b0m_v0m_n263 
  // sz:2: index:4 c0sm_b0m_rdata[0] c0sm_b0m_rdata[1] 
  // sz:2: index:5 c0sm_b0m_v0m_n331 c0sm_b0m_v0m_n332 
  // sz:2: index:6 s0m_m0m_n1 s0m_m0m_n1 
  // sz:2: index:7 s0m_request1[0] s0m_request1[0] 
  // sz:2: index:8 s0m_m0m_n3 s0m_m0m_n2 
  // sz:2: index:9 s0m_m1m_n1 s0m_m1m_n1 
  // sz:2: index:10 s0m_request1[1] s0m_request1[1] 
  // sz:2: index:11 s0m_m1m_n3 s0m_m1m_n2 
  // sz:12: index:12 flitout_switch_0[6] flitout_switch_0[5] flitout_switch_0[4] flitout_switch_0[3] flitout_switch_0[7] flitout_switch_0[8] flitout_switch_0[9] flitout_switch_0[0] flitout_switch_0[10] flitout_switch_0[2] flitout_switch_0[11] flitout_switch_0[1] 
  // sz:12: index:13 flitout_switch_1[6] flitout_switch_1[5] flitout_switch_1[4] flitout_switch_1[3] flitout_switch_1[7] flitout_switch_1[8] flitout_switch_1[9] flitout_switch_1[0] flitout_switch_1[10] flitout_switch_1[2] flitout_switch_1[11] flitout_switch_1[1] 
  // sz:12: index:14 x0m_bx6m_m0m_int01 x0m_bx5m_m0m_int01 x0m_bx4m_m0m_int01 x0m_bx3m_m0m_int01 x0m_bx7m_m0m_int01 x0m_bx8m_m0m_int01 x0m_bx9m_m0m_int01 x0m_bx0m_m0m_int01 x0m_bx10m_m0m_int01 x0m_bx2m_m0m_int01 x0m_bx11m_m0m_int01 x0m_bx1m_m0m_int01 
  // sz:12: index:15 x0m_bx6m_m0m_int01 x0m_bx5m_m0m_int01 x0m_bx4m_m0m_int01 x0m_bx3m_m0m_int01 x0m_bx2m_m0m_int01 x0m_bx1m_m0m_int01 x0m_bx11m_m0m_int01 x0m_bx0m_m0m_int01 x0m_bx10m_m0m_int01 x0m_bx7m_m0m_int01 x0m_bx8m_m0m_int01 x0m_bx9m_m0m_int01 
  // sz:12: index:16 x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic1_ x0m__logic0_ x0m__logic1_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ 
  // sz:12: index:17 flitout_0[6] flitout_0[5] flitout_0[4] flitout_0[3] flitout_0[2] flitout_0[1] flitout_0[11] flitout_0[0] flitout_0[10] flitout_0[7] flitout_0[8] flitout_0[9] 
  // sz:11: index:18 flitout_switch_0[5] flitout_switch_0[4] flitout_switch_0[3] flitout_switch_0[7] flitout_switch_0[2] flitout_switch_0[8] flitout_switch_0[9] flitout_switch_0[0] flitout_switch_0[10] flitout_switch_0[11] flitout_switch_0[1] 
  // sz:11: index:19 flitout_switch_1[5] flitout_switch_1[4] flitout_switch_1[3] flitout_switch_1[7] flitout_switch_1[2] flitout_switch_1[8] flitout_switch_1[9] flitout_switch_1[0] flitout_switch_1[10] flitout_switch_1[11] flitout_switch_1[1] 
  // sz:11: index:20 x0m_bx5m_m1m_int01 x0m_bx4m_m1m_int01 x0m_bx3m_m1m_int01 x0m_bx7m_m1m_int01 x0m_bx2m_m1m_int01 x0m_bx8m_m1m_int01 x0m_bx9m_m1m_int01 x0m_bx0m_m1m_int01 x0m_bx10m_m1m_int01 x0m_bx11m_m1m_int01 x0m_bx1m_m1m_int01 
  // sz:12: index:21 x0m_bx11m_m1m_int01 x0m_bx3m_m1m_int01 x0m_bx1m_m1m_int01 x0m_bx2m_m1m_int01 x0m_bx0m_m1m_int01 x0m_bx10m_m1m_int01 x0m_bx6m_m1m_int01 x0m_bx7m_m1m_int01 x0m_bx8m_m1m_int01 x0m_bx9m_m1m_int01 x0m_bx5m_m1m_int01 x0m_bx4m_m1m_int01 
  // sz:12: index:22 x0m__logic0_ x0m__logic0_ x0m__logic1_ x0m__logic0_ x0m__logic1_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ 
  // sz:12: index:23 flitout_1[11] flitout_1[3] flitout_1[1] flitout_1[2] flitout_1[0] flitout_1[10] flitout_1[6] flitout_1[7] flitout_1[8] flitout_1[9] flitout_1[5] flitout_1[4] 
  // sz:2: index:24 c0nm_b0m_v0m_n105 c0nm_b0m_v0m_n122 
  // sz:2: index:25 c0nm_b0m_v0m_n106 c0nm_b0m_v0m_n123 
  // sz:2: index:26 c0nm_b0m_v0m_n219 c0nm_b0m_v0m_n218 
  // sz:2: index:27 c0nm_b0m_v0m_n61 c0nm_b0m_v0m_n60 
  // sz:2: index:28 c0nm_b0m_v0m_n97 c0nm_b0m_v0m_n101 
  // sz:2: index:29 c0nm_b0m_v0m_n231 c0nm_b0m_v0m_n230 
  // sz:2: index:30 c0nm_b0m_v0m_n74 c0nm_b0m_v0m_n79 
  // sz:2: index:31 c0nm_b0m_v0m_n75 c0nm_b0m_v0m_n80 
  // sz:2: index:32 c0nm_b0m_v0m_n243 c0nm_b0m_v0m_n242 
  // sz:2: index:33 c0nm_b0m_v0m_n23 c0nm_b0m_v0m_n29 
  // sz:2: index:34 c0nm_b0m_v0m_n24 c0nm_b0m_v0m_n30 
  // sz:2: index:35 c0nm_b0m_v0m_n254 c0nm_b0m_v0m_n253 
  // sz:2: index:36 c0nm_v0m_n7 c0nm_v0m_n3 
  // sz:2: index:37 c0nm_routewire[0] c0nm_routewire[1] 
  // sz:2: index:38 c0nm_v0m_n6 c0nm_v0m_n2 
  // sz:2: index:39 c0nm_v0m_state_queuelen_0_ c0nm_v0m_n20 
  // sz:2: index:40 c0nm_v0m_n18 c0nm_v0m_n21 
  // sz:2: index:41 c0nm_v0m_n15 c0nm_v0m_n19 
  // sz:2: index:42 c0sm_b0m_v0m_n105 c0sm_b0m_v0m_n122 
  // sz:2: index:43 c0sm_b0m_v0m_n106 c0sm_b0m_v0m_n123 
  // sz:2: index:44 c0sm_b0m_v0m_n319 c0sm_b0m_v0m_n320 
  // sz:2: index:45 c0sm_b0m_v0m_n344 c0sm_b0m_v0m_n343 
  // sz:2: index:46 c0sm_b0m_v0m_n101 c0sm_b0m_v0m_n97 
  // sz:2: index:47 c0sm_b0m_v0m_n308 c0sm_b0m_v0m_n307 
  // sz:2: index:48 c0sm_b0m_v0m_n79 c0sm_b0m_v0m_n74 
  // sz:2: index:49 c0sm_b0m_v0m_n80 c0sm_b0m_v0m_n75 
  // sz:2: index:50 c0sm_b0m_v0m_n296 c0sm_b0m_v0m_n295 
  // sz:2: index:51 c0sm_b0m_v0m_n29 c0sm_b0m_v0m_n23 
  // sz:2: index:52 c0sm_b0m_v0m_n30 c0sm_b0m_v0m_n24 
  // sz:2: index:53 c0sm_b0m_v0m_n285 c0sm_b0m_v0m_n284 
  // sz:2: index:54 c0sm_v0m_n7 c0sm_v0m_n3 
  // sz:2: index:55 c0sm_routewire[0] c0sm_routewire[1] 
  // sz:2: index:56 c0sm_v0m_n6 c0sm_v0m_n2 
  // sz:2: index:57 c0sm_v0m_state_queuelen_0_ c0sm_v0m_n20 
  // sz:2: index:58 c0sm_v0m_n18 c0sm_v0m_n21 
  // sz:2: index:59 c0sm_v0m_n15 c0sm_v0m_n19 
  // sz:2: index:60 s0m_n13 s0m_n17 
  // sz:2: index:61 s0m_n14 s0m_n18 
  // sz:2: index:62 s0m_n23 s0m_n22 
  // sz:2: index:63 s0m_n6 s0m_n10 
  // sz:2: index:64 s0m_n7 s0m_n11 
  // sz:2: index:65 s0m_n25 s0m_n24 
  // sz:2: index:66 s0m_n4 s0m_n26 
  // sz:2: index:67 s0m_n5 c0nm_v0m_n9 
  // sz:2: index:68 nomorebufs_0 s0m_debit_outvc0 
  // sz:2: index:69 s0m_n1 s0m_n20 
  // sz:2: index:70 s0m_n2 c0nm_v0m_n9 
  // sz:2: index:71 s0m_tail_outvc1 s0m_debit_outvc1 
  // sz:10: index:72 c0nm_b0m_v0m_n200 c0nm_b0m_v0m_n201 c0nm_b0m_v0m_n202 c0nm_b0m_v0m_n199 c0nm_b0m_v0m_n203 c0nm_b0m_v0m_n204 c0nm_b0m_v0m_n205 c0nm_b0m_v0m_n196 c0nm_b0m_v0m_n197 c0nm_b0m_v0m_n198 
  // sz:10: index:73 c0sm_b0m_v0m_n334 c0sm_b0m_v0m_n335 c0sm_b0m_v0m_n336 c0sm_b0m_v0m_n333 c0sm_b0m_v0m_n337 c0sm_b0m_v0m_n338 c0sm_b0m_v0m_n339 c0sm_b0m_v0m_n340 c0sm_b0m_v0m_n341 c0sm_b0m_v0m_n342 
  // sz:2: index:74 c0nm_r0m_n12 c0sm_r0m_n12 
  // sz:2: index:75 c0nm_b0m_v0m_n127 c0nm_b0m_v0m_n118 
  // sz:20: index:76 c0nm_b0m_v0m_n137 c0nm_b0m_v0m_n137 c0nm_b0m_v0m_n143 c0nm_b0m_v0m_n143 c0nm_b0m_v0m_n185 c0nm_b0m_v0m_n185 c0nm_b0m_v0m_n167 c0nm_b0m_v0m_n167 c0nm_b0m_v0m_n173 c0nm_b0m_v0m_n173 c0nm_b0m_v0m_n179 c0nm_b0m_v0m_n179 c0nm_b0m_v0m_n161 c0nm_b0m_v0m_n161 c0nm_b0m_v0m_n155 c0nm_b0m_v0m_n155 c0nm_b0m_v0m_n149 c0nm_b0m_v0m_n149 c0nm_b0m_v0m_n195 c0nm_b0m_v0m_n195 
  // sz:2: index:77 c0nm_b0m_v0m_n137 c0nm_b0m_v0m_n137 
  // sz:2: index:78 c0nm_b0m_v0m_n143 c0nm_b0m_v0m_n143 
  // sz:2: index:79 c0nm_b0m_v0m_n149 c0nm_b0m_v0m_n149 
  // sz:2: index:80 c0nm_b0m_v0m_n155 c0nm_b0m_v0m_n155 
  // sz:2: index:81 c0nm_b0m_v0m_n161 c0nm_b0m_v0m_n161 
  // sz:2: index:82 c0nm_b0m_v0m_n167 c0nm_b0m_v0m_n167 
  // sz:2: index:83 c0nm_b0m_v0m_n173 c0nm_b0m_v0m_n173 
  // sz:2: index:84 c0nm_b0m_v0m_n179 c0nm_b0m_v0m_n179 
  // sz:2: index:85 c0nm_b0m_v0m_n185 c0nm_b0m_v0m_n185 
  // sz:2: index:86 c0nm_b0m_v0m_n195 c0nm_b0m_v0m_n195 
  // sz:12: index:87 c0nm_b0m_v0m_n269 c0nm_b0m_v0m_n265 c0nm_b0m_v0m_n266 c0nm_b0m_v0m_n267 c0nm_b0m_v0m_n268 c0nm_b0m_v0m_n276 c0nm_b0m_v0m_n270 c0nm_b0m_v0m_n275 c0nm_b0m_v0m_n274 c0nm_b0m_v0m_n273 c0nm_b0m_v0m_n272 c0nm_b0m_v0m_n271 
  // sz:2: index:88 c0nm_b0m_v0m_n274 c0nm_b0m_v0m_n182 
  // sz:2: index:89 c0nm_b0m_v0m_n273 c0nm_b0m_v0m_n189 
  // sz:2: index:90 c0nm_b0m_v0m_n272 c0nm_b0m_v0m_n133 
  // sz:2: index:91 c0nm_b0m_v0m_n271 c0nm_b0m_v0m_n140 
  // sz:2: index:92 c0nm_b0m_v0m_n270 c0nm_b0m_v0m_n146 
  // sz:2: index:93 c0nm_b0m_v0m_n269 c0nm_b0m_v0m_n152 
  // sz:2: index:94 c0nm_b0m_v0m_n268 c0nm_b0m_v0m_n158 
  // sz:2: index:95 c0nm_b0m_v0m_n267 c0nm_b0m_v0m_n164 
  // sz:2: index:96 c0nm_b0m_v0m_n266 c0nm_b0m_v0m_n170 
  // sz:2: index:97 c0nm_b0m_v0m_n265 c0nm_b0m_v0m_n176 
  // sz:12: index:98 c0nm_b0m_v0m_n172 c0nm_b0m_v0m_n126 c0nm_b0m_v0m_n178 c0nm_b0m_v0m_n184 c0nm_b0m_v0m_n117 c0nm_b0m_v0m_n194 c0nm_b0m_v0m_n154 c0nm_b0m_v0m_n160 c0nm_b0m_v0m_n142 c0nm_b0m_v0m_n166 c0nm_b0m_v0m_n136 c0nm_b0m_v0m_n148 
  // sz:10: index:99 c0nm_b0m_v0m_n170 c0nm_b0m_v0m_n146 c0nm_b0m_v0m_n133 c0nm_b0m_v0m_n140 c0nm_b0m_v0m_n152 c0nm_b0m_v0m_n164 c0nm_b0m_v0m_n158 c0nm_b0m_v0m_n189 c0nm_b0m_v0m_n182 c0nm_b0m_v0m_n176 
  // sz:2: index:100 c0sm_b0m_v0m_n127 c0sm_b0m_v0m_n118 
  // sz:20: index:101 c0sm_b0m_v0m_n143 c0sm_b0m_v0m_n143 c0sm_b0m_v0m_n137 c0sm_b0m_v0m_n137 c0sm_b0m_v0m_n149 c0sm_b0m_v0m_n149 c0sm_b0m_v0m_n195 c0sm_b0m_v0m_n195 c0sm_b0m_v0m_n185 c0sm_b0m_v0m_n185 c0sm_b0m_v0m_n179 c0sm_b0m_v0m_n179 c0sm_b0m_v0m_n173 c0sm_b0m_v0m_n173 c0sm_b0m_v0m_n167 c0sm_b0m_v0m_n167 c0sm_b0m_v0m_n161 c0sm_b0m_v0m_n161 c0sm_b0m_v0m_n155 c0sm_b0m_v0m_n155 
  // sz:2: index:102 c0sm_b0m_v0m_n137 c0sm_b0m_v0m_n137 
  // sz:2: index:103 c0sm_b0m_v0m_n143 c0sm_b0m_v0m_n143 
  // sz:2: index:104 c0sm_b0m_v0m_n149 c0sm_b0m_v0m_n149 
  // sz:2: index:105 c0sm_b0m_v0m_n155 c0sm_b0m_v0m_n155 
  // sz:2: index:106 c0sm_b0m_v0m_n161 c0sm_b0m_v0m_n161 
  // sz:2: index:107 c0sm_b0m_v0m_n167 c0sm_b0m_v0m_n167 
  // sz:2: index:108 c0sm_b0m_v0m_n173 c0sm_b0m_v0m_n173 
  // sz:2: index:109 c0sm_b0m_v0m_n179 c0sm_b0m_v0m_n179 
  // sz:2: index:110 c0sm_b0m_v0m_n185 c0sm_b0m_v0m_n185 
  // sz:2: index:111 c0sm_b0m_v0m_n195 c0sm_b0m_v0m_n195 
  // sz:12: index:112 c0sm_b0m_v0m_n272 c0sm_b0m_v0m_n273 c0sm_b0m_v0m_n274 c0sm_b0m_v0m_n271 c0sm_b0m_v0m_n270 c0sm_b0m_v0m_n275 c0sm_b0m_v0m_n269 c0sm_b0m_v0m_n268 c0sm_b0m_v0m_n267 c0sm_b0m_v0m_n276 c0sm_b0m_v0m_n265 c0sm_b0m_v0m_n266 
  // sz:2: index:113 c0sm_b0m_v0m_n274 c0sm_b0m_v0m_n182 
  // sz:2: index:114 c0sm_b0m_v0m_n273 c0sm_b0m_v0m_n189 
  // sz:2: index:115 c0sm_b0m_v0m_n272 c0sm_b0m_v0m_n133 
  // sz:2: index:116 c0sm_b0m_v0m_n271 c0sm_b0m_v0m_n140 
  // sz:2: index:117 c0sm_b0m_v0m_n270 c0sm_b0m_v0m_n146 
  // sz:2: index:118 c0sm_b0m_v0m_n269 c0sm_b0m_v0m_n152 
  // sz:2: index:119 c0sm_b0m_v0m_n268 c0sm_b0m_v0m_n158 
  // sz:2: index:120 c0sm_b0m_v0m_n267 c0sm_b0m_v0m_n164 
  // sz:2: index:121 c0sm_b0m_v0m_n266 c0sm_b0m_v0m_n170 
  // sz:2: index:122 c0sm_b0m_v0m_n265 c0sm_b0m_v0m_n176 
  // sz:12: index:123 c0sm_b0m_v0m_n184 c0sm_b0m_v0m_n194 c0sm_b0m_v0m_n142 c0sm_b0m_v0m_n136 c0sm_b0m_v0m_n126 c0sm_b0m_v0m_n117 c0sm_b0m_v0m_n178 c0sm_b0m_v0m_n172 c0sm_b0m_v0m_n166 c0sm_b0m_v0m_n160 c0sm_b0m_v0m_n154 c0sm_b0m_v0m_n148 
  // sz:10: index:124 c0sm_b0m_v0m_n170 c0sm_b0m_v0m_n133 c0sm_b0m_v0m_n164 c0sm_b0m_v0m_n140 c0sm_b0m_v0m_n158 c0sm_b0m_v0m_n146 c0sm_b0m_v0m_n152 c0sm_b0m_v0m_n189 c0sm_b0m_v0m_n182 c0sm_b0m_v0m_n176 
  // sz:12: index:125 flitout_switch_0[6] flitout_switch_0[5] flitout_switch_0[4] flitout_switch_0[3] flitout_switch_0[2] flitout_switch_0[1] flitout_switch_0[11] flitout_switch_0[0] flitout_switch_0[10] flitout_switch_0[7] flitout_switch_0[8] flitout_switch_0[9] 
  // sz:12: index:126 flitout_switch_1[6] flitout_switch_1[5] flitout_switch_1[4] flitout_switch_1[3] flitout_switch_1[2] flitout_switch_1[1] flitout_switch_1[11] flitout_switch_1[0] flitout_switch_1[10] flitout_switch_1[7] flitout_switch_1[8] flitout_switch_1[9] 
  // sz:11: index:127 flitout_switch_0[3] flitout_switch_0[1] flitout_switch_0[2] flitout_switch_0[0] flitout_switch_0[10] flitout_switch_0[6] flitout_switch_0[7] flitout_switch_0[8] flitout_switch_0[9] flitout_switch_0[5] flitout_switch_0[4] 
  // sz:11: index:128 flitout_switch_1[3] flitout_switch_1[1] flitout_switch_1[2] flitout_switch_1[0] flitout_switch_1[10] flitout_switch_1[6] flitout_switch_1[7] flitout_switch_1[8] flitout_switch_1[9] flitout_switch_1[5] flitout_switch_1[4] 
  // sz:11: index:129 x0m__logic0_ x0m__logic1_ x0m__logic0_ x0m__logic1_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ 
  // sz:11: index:130 flitout_1[3] flitout_1[1] flitout_1[2] flitout_1[0] flitout_1[10] flitout_1[6] flitout_1[7] flitout_1[8] flitout_1[9] flitout_1[5] flitout_1[4] 
  // sz:10: index:131 c0nm_b0m_v0m_n208 c0nm_b0m_v0m_n209 c0nm_b0m_v0m_n210 c0nm_b0m_v0m_n211 c0nm_b0m_v0m_n212 c0nm_b0m_v0m_n213 c0nm_b0m_v0m_n214 c0nm_b0m_v0m_n215 c0nm_b0m_v0m_n216 c0nm_b0m_v0m_n217 
  // sz:10: index:132 c0nm_b0m_v0m_n222 c0nm_b0m_v0m_n229 c0nm_b0m_v0m_n228 c0nm_b0m_v0m_n227 c0nm_b0m_v0m_n226 c0nm_b0m_v0m_n225 c0nm_b0m_v0m_n224 c0nm_b0m_v0m_n223 c0nm_b0m_v0m_n221 c0nm_b0m_v0m_n220 
  // sz:10: index:133 c0nm_b0m_v0m_n232 c0nm_b0m_v0m_n239 c0nm_b0m_v0m_n238 c0nm_b0m_v0m_n237 c0nm_b0m_v0m_n236 c0nm_b0m_v0m_n235 c0nm_b0m_v0m_n234 c0nm_b0m_v0m_n233 c0nm_b0m_v0m_n241 c0nm_b0m_v0m_n240 
  // sz:10: index:134 c0nm_b0m_v0m_n247 c0nm_b0m_v0m_n255 c0nm_b0m_v0m_n252 c0nm_b0m_v0m_n251 c0nm_b0m_v0m_n250 c0nm_b0m_v0m_n249 c0nm_b0m_v0m_n248 c0nm_b0m_v0m_n246 c0nm_b0m_v0m_n245 c0nm_b0m_v0m_n244 
  // sz:10: index:135 c0sm_b0m_v0m_n321 c0sm_b0m_v0m_n322 c0sm_b0m_v0m_n323 c0sm_b0m_v0m_n324 c0sm_b0m_v0m_n325 c0sm_b0m_v0m_n326 c0sm_b0m_v0m_n327 c0sm_b0m_v0m_n328 c0sm_b0m_v0m_n329 c0sm_b0m_v0m_n330 
  // sz:10: index:136 c0sm_b0m_v0m_n309 c0sm_b0m_v0m_n310 c0sm_b0m_v0m_n311 c0sm_b0m_v0m_n312 c0sm_b0m_v0m_n313 c0sm_b0m_v0m_n314 c0sm_b0m_v0m_n315 c0sm_b0m_v0m_n316 c0sm_b0m_v0m_n317 c0sm_b0m_v0m_n318 
  // sz:10: index:137 c0sm_b0m_v0m_n301 c0sm_b0m_v0m_n300 c0sm_b0m_v0m_n299 c0sm_b0m_v0m_n298 c0sm_b0m_v0m_n297 c0sm_b0m_v0m_n302 c0sm_b0m_v0m_n305 c0sm_b0m_v0m_n306 c0sm_b0m_v0m_n304 c0sm_b0m_v0m_n303 
  // sz:10: index:138 c0sm_b0m_v0m_n288 c0sm_b0m_v0m_n294 c0sm_b0m_v0m_n293 c0sm_b0m_v0m_n292 c0sm_b0m_v0m_n291 c0sm_b0m_v0m_n290 c0sm_b0m_v0m_n289 c0sm_b0m_v0m_n287 c0sm_b0m_v0m_n286 c0sm_b0m_v0m_n283 
  // sz:2: index:139 c0sm_r0m_n7 c0nm_r0m_n7 
  // sz:4: index:140 c0nm_b0m_v0m_n80 c0nm_b0m_v0m_n101 c0nm_b0m_v0m_n30 c0nm_b0m_v0m_n123 
  // sz:4: index:141 c0nm_b0m_v0m_n24 c0nm_b0m_v0m_n106 c0nm_b0m_v0m_n75 c0nm_b0m_v0m_n97 
  // sz:2: index:142 c0nm_b0m_v0m_n101 c0nm_b0m_v0m_n97 
  // sz:2: index:143 c0nm_b0m_v0m_n80 c0nm_b0m_v0m_n75 
  // sz:4: index:144 c0sm_b0m_v0m_n101 c0sm_b0m_v0m_n123 c0sm_b0m_v0m_n80 c0sm_b0m_v0m_n30 
  // sz:4: index:145 c0sm_b0m_v0m_n106 c0sm_b0m_v0m_n97 c0sm_b0m_v0m_n75 c0sm_b0m_v0m_n24 
  // sz:2: index:146 c0nm_b0m_v0m_n112 c0nm_b0m_v0m_n124 
  // sz:2: index:147 c0nm_b0m_v0m_n112 c0nm_b0m_v0m_n112 
  // sz:2: index:148 c0nm_b0m_v0m_n124 c0nm_b0m_v0m_n124 
  // sz:4: index:149 c0nm_b0m_v0m_n112 c0nm_b0m_v0m_n112 c0nm_b0m_v0m_n124 c0nm_b0m_v0m_n124 
  // sz:4: index:150 c0nm_b0m_v0m_n112 c0nm_b0m_v0m_n112 c0nm_b0m_v0m_n112 c0nm_b0m_v0m_n112 
  // sz:4: index:151 c0nm_b0m_v0m_n124 c0nm_b0m_v0m_n124 c0nm_b0m_v0m_n124 c0nm_b0m_v0m_n124 
  // sz:2: index:152 c0sm_b0m_v0m_n112 c0sm_b0m_v0m_n124 
  // sz:2: index:153 c0sm_b0m_v0m_n112 c0sm_b0m_v0m_n112 
  // sz:2: index:154 c0sm_b0m_v0m_n124 c0sm_b0m_v0m_n124 
  // sz:4: index:155 c0sm_b0m_v0m_n112 c0sm_b0m_v0m_n112 c0sm_b0m_v0m_n124 c0sm_b0m_v0m_n124 
  // sz:4: index:156 c0sm_b0m_v0m_n112 c0sm_b0m_v0m_n112 c0sm_b0m_v0m_n112 c0sm_b0m_v0m_n112 
  // sz:4: index:157 c0sm_b0m_v0m_n124 c0sm_b0m_v0m_n124 c0sm_b0m_v0m_n124 c0sm_b0m_v0m_n124 
  // sz:4: index:158 c0nm_b0m_v0m_n264 c0nm_r0m_n14 c0nm_r0m_n8 c0nm_r0m_n9 
  // sz:2: index:159 c0nm_r0m_n14 c0nm_b0m_v0m_n36 
  // sz:2: index:160 c0nm_r0m_n9 c0nm_b0m_v0m_n42 
  // sz:2: index:161 c0nm_r0m_n8 c0nm_b0m_v0m_n45 
  // sz:10: index:162 c0nm_b0m_v0m_n33 c0nm_b0m_v0m_n36 c0nm_b0m_v0m_n69 c0nm_b0m_v0m_n66 c0nm_b0m_v0m_n39 c0nm_b0m_v0m_n42 c0nm_b0m_v0m_n63 c0nm_b0m_v0m_n48 c0nm_b0m_v0m_n45 c0nm_b0m_v0m_n17 
  // sz:4: index:163 c0sm_r0m_n14 c0sm_r0m_n9 c0sm_r0m_n8 c0sm_b0m_v0m_n264 
  // sz:2: index:164 c0sm_r0m_n14 c0sm_b0m_v0m_n36 
  // sz:2: index:165 c0sm_r0m_n9 c0sm_b0m_v0m_n42 
  // sz:2: index:166 c0sm_r0m_n8 c0sm_b0m_v0m_n45 
  // sz:10: index:167 c0sm_b0m_v0m_n33 c0sm_b0m_v0m_n48 c0sm_b0m_v0m_n17 c0sm_b0m_v0m_n45 c0sm_b0m_v0m_n42 c0sm_b0m_v0m_n63 c0sm_b0m_v0m_n66 c0sm_b0m_v0m_n39 c0sm_b0m_v0m_n69 c0sm_b0m_v0m_n36 
  // sz:12: index:168 c0nm_headflit[2] c0nm_headflit[0] c0nm_headflit[1] c0nm_headflit[3] c0nm_headflit[4] c0nm_headflit[5] c0nm_headflit[6] c0nm_headflit[7] c0nm_b0m_headflit_9_ c0nm_b0m_headflit_8_ c0nm_b0m_headflit_11_ c0nm_b0m_headflit_10_ 
  // sz:2: index:169 c0nm_headflit[0] c0nm_b0m_v0m_n27 
  // sz:2: index:170 c0nm_headflit[1] c0nm_b0m_v0m_n32 
  // sz:2: index:171 c0nm_b0m_headflit_10_ c0nm_b0m_v0m_n181 
  // sz:2: index:172 c0nm_b0m_headflit_11_ c0nm_b0m_v0m_n188 
  // sz:2: index:173 c0nm_headflit[2] c0nm_b0m_v0m_n132 
  // sz:2: index:174 c0nm_headflit[3] c0nm_b0m_v0m_n139 
  // sz:2: index:175 c0nm_headflit[4] c0nm_b0m_v0m_n145 
  // sz:2: index:176 c0nm_headflit[5] c0nm_b0m_v0m_n151 
  // sz:2: index:177 c0nm_headflit[6] c0nm_b0m_v0m_n157 
  // sz:2: index:178 c0nm_headflit[7] c0nm_b0m_v0m_n163 
  // sz:2: index:179 c0nm_b0m_headflit_8_ c0nm_b0m_v0m_n169 
  // sz:2: index:180 c0nm_b0m_headflit_9_ c0nm_b0m_v0m_n175 
  // sz:12: index:181 c0nm_b0m_v0m_n139 c0nm_b0m_v0m_n132 c0nm_b0m_v0m_n145 c0nm_b0m_v0m_n169 c0nm_b0m_v0m_n188 c0nm_b0m_v0m_n181 c0nm_b0m_v0m_n175 c0nm_b0m_v0m_n163 c0nm_b0m_v0m_n157 c0nm_b0m_v0m_n151 c0nm_b0m_v0m_n27 c0nm_b0m_v0m_n32 
  // sz:12: index:182 c0sm_headflit[5] c0sm_headflit[0] c0sm_headflit[1] c0sm_headflit[2] c0sm_headflit[3] c0sm_headflit[4] c0sm_headflit[6] c0sm_headflit[7] c0sm_b0m_headflit_11_ c0sm_b0m_headflit_10_ c0sm_b0m_headflit_8_ c0sm_b0m_headflit_9_ 
  // sz:2: index:183 c0sm_headflit[0] c0sm_b0m_v0m_n27 
  // sz:2: index:184 c0sm_headflit[1] c0sm_b0m_v0m_n32 
  // sz:2: index:185 c0sm_b0m_headflit_10_ c0sm_b0m_v0m_n181 
  // sz:2: index:186 c0sm_b0m_headflit_11_ c0sm_b0m_v0m_n188 
  // sz:2: index:187 c0sm_headflit[2] c0sm_b0m_v0m_n132 
  // sz:2: index:188 c0sm_headflit[3] c0sm_b0m_v0m_n139 
  // sz:2: index:189 c0sm_headflit[4] c0sm_b0m_v0m_n145 
  // sz:2: index:190 c0sm_headflit[5] c0sm_b0m_v0m_n151 
  // sz:2: index:191 c0sm_headflit[6] c0sm_b0m_v0m_n157 
  // sz:2: index:192 c0sm_headflit[7] c0sm_b0m_v0m_n163 
  // sz:2: index:193 c0sm_b0m_headflit_8_ c0sm_b0m_v0m_n169 
  // sz:2: index:194 c0sm_b0m_headflit_9_ c0sm_b0m_v0m_n175 
  // sz:12: index:195 c0sm_b0m_v0m_n32 c0sm_b0m_v0m_n151 c0sm_b0m_v0m_n157 c0sm_b0m_v0m_n145 c0sm_b0m_v0m_n175 c0sm_b0m_v0m_n181 c0sm_b0m_v0m_n169 c0sm_b0m_v0m_n188 c0sm_b0m_v0m_n163 c0sm_b0m_v0m_n27 c0sm_b0m_v0m_n139 c0sm_b0m_v0m_n132 
  // sz:2: index:196 c0sm_r0m_n16 c0nm_r0m_n16 
  // sz:10: index:197 c0nm_b0m_wdata_11_ c0nm_b0m_wdata_8_ c0nm_b0m_wdata_9_ c0nm_b0m_wdata_7_ c0nm_b0m_wdata_6_ c0nm_b0m_wdata_5_ c0nm_b0m_wdata_4_ c0nm_b0m_wdata_3_ c0nm_b0m_wdata_2_ c0nm_b0m_wdata_10_ 
  // sz:10: index:198 flitout_switch_0[11] flitout_switch_0[6] flitout_switch_0[5] flitout_switch_0[4] flitout_switch_0[3] flitout_switch_0[2] flitout_switch_0[10] flitout_switch_0[9] flitout_switch_0[8] flitout_switch_0[7] 
  // sz:2: index:199 c0nm_b0m_v0m_n115 c0nm_b0m_v0m_n113 
  // sz:2: index:200 s0m_request0[1] c0nm_v0m_n3 
  // sz:2: index:201 s0m_request0[0] c0nm_v0m_n7 
  // sz:10: index:202 c0sm_b0m_wdata_10_ c0sm_b0m_wdata_9_ c0sm_b0m_wdata_8_ c0sm_b0m_wdata_7_ c0sm_b0m_wdata_6_ c0sm_b0m_wdata_5_ c0sm_b0m_wdata_4_ c0sm_b0m_wdata_3_ c0sm_b0m_wdata_11_ c0sm_b0m_wdata_2_ 
  // sz:10: index:203 flitout_switch_1[5] flitout_switch_1[9] flitout_switch_1[8] flitout_switch_1[7] flitout_switch_1[6] flitout_switch_1[4] flitout_switch_1[3] flitout_switch_1[2] flitout_switch_1[11] flitout_switch_1[10] 
  // sz:2: index:204 c0sm_v0m_n3 c0sm_v0m_n7 
  // sz:2: index:205 c0sm_b0m_v0m_n113 c0sm_b0m_v0m_n115 
  // sz:2: index:206 s0m_request1[1] c0sm_v0m_n3 
  // sz:2: index:207 s0m_request1[0] c0sm_v0m_n7 
  // sz:2: index:208 s0m_request0[0] s0m_request1[0] 
  // sz:2: index:209 s0m_request0[1] s0m_request1[1] 
  // sz:2: index:210 c0nm_r0m_n15 c0sm_r0m_n15 
  // sz:20: index:211 x0m_n3 x0m_n4 x0m_n5 x0m_n6 c0nm_v0m_n1 c0sm_v0m_n1 c0sm_b0m_v0m_n1 c0nm_b0m_v0m_n1 c0sm_b0m_v0m_n81 c0sm_b0m_v0m_n2 c0sm_b0m_v0m_n129 c0sm_b0m_v0m_n102 c0nm_b0m_v0m_n2 c0nm_b0m_v0m_n81 c0nm_b0m_v0m_n102 c0nm_b0m_v0m_n129 c0sm_b0m_v0m_n262 c0nm_b0m_v0m_n262 c0nm_b0m_v0m_n263 c0sm_b0m_v0m_n263 
  // sz:3: index:212 c0nm_b0m_v0m_n1 c0nm_b0m_v0m_n135 c0nm_b0m_v0m_n116 
  // sz:2: index:213 c0nm_b0m_v0m_n102 c0nm_b0m_v0m_n135 
  // sz:3: index:214 c0sm_b0m_v0m_n1 c0sm_b0m_v0m_n135 c0sm_b0m_v0m_n116 
  // sz:2: index:215 c0sm_b0m_v0m_n135 c0sm_b0m_v0m_n102 
  // sz:2: index:216 flitout_0[1] flitout_0[0] 
  // sz:2: index:217 flitout_1[1] flitout_1[0] 
  // sz:2: index:218 c0nm_n2 c0nm_b0m_n1 
  // sz:2: index:219 c0sm_n3 c0sm_b0m_n2 
  // sz:14: index:220 c0sm_b0m_v0m_n20 c0nm_b0m_v0m_n20 c0sm_b0m_v0m_n81 c0sm_b0m_v0m_n2 c0sm_b0m_v0m_n129 c0sm_b0m_v0m_n102 c0nm_b0m_v0m_n2 c0nm_b0m_v0m_n81 c0nm_b0m_v0m_n102 c0nm_b0m_v0m_n129 c0nm_b0m_v0m_n263 c0sm_b0m_v0m_n263 s0m_o0nm_n36 s0m_o0sm_n36 
  // sz:2: index:221 s0m_n3 s0m_n1 
  // sz:2: index:222 s0m_n26 s0m_n20 
  // sz:2: index:223 s0m_n18 s0m_n14 
  // sz:2: index:224 s0m_n11 s0m_n7 
  // sz:2: index:225 s0m_n3 s0m_n26 
  // sz:30: index:226 c0sm_v0m_n8 c0nm_v0m_n8 s0m_n9 s0m_n16 c0nm_b0m_v0m_n8 c0sm_b0m_v0m_n8 s0m_o0nm_n3 s0m_o0sm_n3 s0m_m0m_n10 s0m_m0m_n10 c0nm_b0m_n9 c0nm_b0m_v0m_n11 c0sm_b0m_v0m_n11 s0m_m1m_n10 s0m_m1m_n10 c0sm_b0m_n9 creditout_0 creditout_1 c0sm_b0m_v0m_n10 c0sm_b0m_v0m_n10 c0nm_b0m_v0m_n10 c0nm_b0m_v0m_n10 c0sm_v0m_n64 c0nm_v0m_n64 c0sm_v0m_n61 c0nm_v0m_n61 c0sm_v0m_n62 c0nm_v0m_n62 s0m_o0nm_n38 s0m_o0sm_n38 
  // sz:5: index:227 c0nm_b0m_v0m_n8 c0nm_b0m_v0m_n119 c0nm_b0m_v0m_n120 c0nm_b0m_v0m_n121 c0nm_b0m_v0m_n128 
  // sz:2: index:228 c0nm_v0m_n8 s0m_n9 
  // sz:4: index:229 c0nm_v0m_n13 c0nm_b0m_n9 creditout_0 c0nm_b0m_v0m_n10 
  // sz:3: index:230 c0nm_b0m_v0m_n115 c0nm_b0m_v0m_n113 c0nm_b0m_v0m_n11 
  // sz:2: index:231 c0nm_v0m_n31 c0nm_v0m_n30 
  // sz:5: index:232 c0sm_b0m_v0m_n8 c0sm_b0m_v0m_n119 c0sm_b0m_v0m_n120 c0sm_b0m_v0m_n121 c0sm_b0m_v0m_n128 
  // sz:2: index:233 c0sm_v0m_n8 s0m_n16 
  // sz:4: index:234 c0sm_v0m_n13 c0sm_b0m_n9 creditout_1 c0sm_b0m_v0m_n10 
  // sz:3: index:235 c0sm_b0m_v0m_n11 c0sm_b0m_v0m_n113 c0sm_b0m_v0m_n115 
  // sz:2: index:236 c0sm_v0m_n32 c0sm_v0m_n33 
  // sz:2: index:237 s0m_m0m_n2 s0m_m1m_n2 
  // sz:4: index:238 x0m_bx4m_m1m_int01 x0m_bx0m_m1m_int01 x0m_bx11m_m1m_int01 x0m_bx1m_m1m_int01 
  // sz:2: index:239 flitout_1[11] flitout_1[4] 
  // sz:5: index:240 c0nm_b0m_v0m_n269 c0nm_b0m_v0m_n268 c0nm_b0m_v0m_n276 c0nm_b0m_v0m_n275 c0nm_b0m_v0m_n271 
  // sz:3: index:241 c0sm_b0m_v0m_n271 c0sm_b0m_v0m_n269 c0sm_b0m_v0m_n268 
  // sz:8: index:242 flitout_1[3] flitout_1[2] flitout_1[10] flitout_1[6] flitout_1[7] flitout_1[8] flitout_1[9] flitout_1[5] 
  // sz:3: index:243 c0nm_r0m_n14 c0nm_r0m_n8 c0nm_r0m_n9 
  // sz:3: index:244 c0sm_r0m_n14 c0sm_r0m_n9 c0sm_r0m_n8 
  // sz:2: index:245 c0sm_b0m_v0m_n32 c0sm_b0m_v0m_n27 
  // sz:2: index:246 c0nm_b0m_v0m_n135 c0nm_b0m_v0m_n116 
  // sz:2: index:247 c0sm_b0m_v0m_n135 c0sm_b0m_v0m_n116 
  // sz:4: index:248 c0sm_b0m_v0m_n20 c0nm_b0m_v0m_n20 s0m_o0nm_n36 s0m_o0sm_n36 
  // sz:26: index:249 s0m_n9 s0m_n16 c0nm_b0m_v0m_n8 c0sm_b0m_v0m_n8 s0m_o0nm_n3 s0m_o0sm_n3 s0m_m0m_n10 s0m_m0m_n10 c0nm_b0m_v0m_n11 c0sm_b0m_v0m_n11 s0m_m1m_n10 s0m_m1m_n10 creditout_0 creditout_1 c0sm_b0m_v0m_n10 c0sm_b0m_v0m_n10 c0nm_b0m_v0m_n10 c0nm_b0m_v0m_n10 c0sm_v0m_n64 c0nm_v0m_n64 c0sm_v0m_n61 c0nm_v0m_n61 c0sm_v0m_n62 c0nm_v0m_n62 s0m_o0nm_n38 s0m_o0sm_n38 
  // sz:2: index:250 c0nm_b0m_v0m_n120 c0nm_b0m_v0m_n121 
  // sz:2: index:251 c0nm_v0m_n13 c0nm_b0m_n9 
  // sz:2: index:252 c0sm_b0m_v0m_n120 c0sm_b0m_v0m_n121 
  // sz:2: index:253 c0sm_v0m_n13 c0sm_b0m_n9 
  // BSIM@ modules: mx245 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx406 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx406 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx248 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx248 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx407 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx407 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx245 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx404 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx404 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx247 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx247 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx405 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx405 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx246 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx246 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   TIELO_X1M_A12TR c0nm_u2 (.Y(c0nm__logic0_));
  TIELO_X1M_A12TR c0nm_b0m_u3 (.Y(c0nm_b0m__logic0_));
  DFFQ_X1M_A12TR c0nm_b0m_dqenablereg_reg (.CK(clk), .Q(c0nm_b0m_dqenablereg), .D(c0nm_b0m_n9));
  // BSIM@ modules: mx374 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u255 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n180), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n71), .C0(c0nm_b0m_v0m_n274), .Y(c0nm_b0m_headflit_10_));
  // BSIM@ modules: mx374 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u250 (.A0(c0nm_b0m_v0m_n186), .A1(c0nm_b0m_v0m_n187), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n21), .C0(c0nm_b0m_v0m_n273), .Y(c0nm_b0m_headflit_11_));
  // BSIM@ modules: mx374 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u215 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n168), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n65), .C0(c0nm_b0m_v0m_n266), .Y(c0nm_b0m_headflit_8_));
  // BSIM@ modules: mx374 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u210 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n174), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n68), .C0(c0nm_b0m_v0m_n265), .Y(c0nm_b0m_headflit_9_));
  // BSIM@ modules: mx343 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR c0nm_b0m_u14 (.A(flitin_0[1]), .B(flitin_0[0]), .Y(c0nm_b0m_n1));
  // BSIM@ modules: mx356 
  // BSIM@ covered_modules=1 :   NOR2B_X0P5M_A12TR c0nm_b0m_u27 (.AN(debitout_0), .B(reset), .Y(c0nm_b0m_n9));
  // BSIM@ modules: mx245 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_0_ (.CK(clk), .Q(c0nm_b0m_rdata[0]), .D(c0nm_b0m_v0m_n207));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_10_ (.CK(clk), .Q(c0nm_b0m_rdata[10]), .D(c0nm_b0m_v0m_n197));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_11_ (.CK(clk), .Q(c0nm_b0m_rdata[11]), .D(c0nm_b0m_v0m_n196));
  // BSIM@ modules: mx245 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_1_ (.CK(clk), .Q(c0nm_b0m_rdata[1]), .D(c0nm_b0m_v0m_n206));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_2_ (.CK(clk), .Q(c0nm_b0m_rdata[2]), .D(c0nm_b0m_v0m_n205));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_3_ (.CK(clk), .Q(c0nm_b0m_rdata[3]), .D(c0nm_b0m_v0m_n204));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_4_ (.CK(clk), .Q(c0nm_b0m_rdata[4]), .D(c0nm_b0m_v0m_n203));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_5_ (.CK(clk), .Q(c0nm_b0m_rdata[5]), .D(c0nm_b0m_v0m_n202));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_6_ (.CK(clk), .Q(c0nm_b0m_rdata[6]), .D(c0nm_b0m_v0m_n201));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_7_ (.CK(clk), .Q(c0nm_b0m_rdata[7]), .D(c0nm_b0m_v0m_n200));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_8_ (.CK(clk), .Q(c0nm_b0m_rdata[8]), .D(c0nm_b0m_v0m_n199));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_9_ (.CK(clk), .Q(c0nm_b0m_rdata[9]), .D(c0nm_b0m_v0m_n198));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_0_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers0_0_), .D(c0nm_b0m_v0m_n243));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_10_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers0_10_), .D(c0nm_b0m_v0m_n233));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_11_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers0_11_), .D(c0nm_b0m_v0m_n232));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_1_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers0_1_), .D(c0nm_b0m_v0m_n242));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_2_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers0_2_), .D(c0nm_b0m_v0m_n241));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_3_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers0_3_), .D(c0nm_b0m_v0m_n240));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_4_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers0_4_), .D(c0nm_b0m_v0m_n239));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_5_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers0_5_), .D(c0nm_b0m_v0m_n238));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_6_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers0_6_), .D(c0nm_b0m_v0m_n237));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_7_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers0_7_), .D(c0nm_b0m_v0m_n236));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_8_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers0_8_), .D(c0nm_b0m_v0m_n235));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers0_reg_9_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers0_9_), .D(c0nm_b0m_v0m_n234));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_0_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers2_0_), .D(c0nm_b0m_v0m_n219));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_10_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers2_10_), .D(c0nm_b0m_v0m_n209));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_11_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers2_11_), .D(c0nm_b0m_v0m_n208));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_1_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers2_1_), .D(c0nm_b0m_v0m_n218));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_2_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers2_2_), .D(c0nm_b0m_v0m_n217));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_3_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers2_3_), .D(c0nm_b0m_v0m_n216));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_4_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers2_4_), .D(c0nm_b0m_v0m_n215));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_5_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers2_5_), .D(c0nm_b0m_v0m_n214));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_6_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers2_6_), .D(c0nm_b0m_v0m_n213));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_7_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers2_7_), .D(c0nm_b0m_v0m_n212));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_8_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers2_8_), .D(c0nm_b0m_v0m_n211));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers2_reg_9_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers2_9_), .D(c0nm_b0m_v0m_n210));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_0_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers3_0_), .D(c0nm_b0m_v0m_n254));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_10_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers3_10_), .D(c0nm_b0m_v0m_n244));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_11_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers3_11_), .D(c0nm_b0m_v0m_n255));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_1_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers3_1_), .D(c0nm_b0m_v0m_n253));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_2_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers3_2_), .D(c0nm_b0m_v0m_n252));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_3_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers3_3_), .D(c0nm_b0m_v0m_n251));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_4_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers3_4_), .D(c0nm_b0m_v0m_n250));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_5_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers3_5_), .D(c0nm_b0m_v0m_n249));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_6_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers3_6_), .D(c0nm_b0m_v0m_n248));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_7_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers3_7_), .D(c0nm_b0m_v0m_n247));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_8_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers3_8_), .D(c0nm_b0m_v0m_n246));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_buffers3_reg_9_ (.CK(clk), .Q(c0nm_b0m_v0m_buffers3_9_), .D(c0nm_b0m_v0m_n245));
  // BSIM@ modules: mx404 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0nm_b0m_v0m_head_reg_0_ (.CK(clk), .Q(c0nm_b0m_v0m_head_0_), .D(c0nm_b0m_v0m_n258));
  // BSIM@ modules: mx404 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0nm_b0m_v0m_head_reg_1_ (.CK(clk), .Q(c0nm_b0m_v0m_head_1_), .D(c0nm_b0m_v0m_n257));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_head_reg_2_ (.CK(clk), .Q(c0nm_b0m_v0m_head_2_), .D(c0nm_b0m_v0m_n256));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u7 (.A(c0nm_b0m_v0m_n8), .Y(c0nm_b0m_v0m_n1));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0nm_b0m_v0m_u208 (.A(c0nm_b0m_v0m_n11), .B(reset), .Y(c0nm_b0m_v0m_n10));
  // BSIM@ modules: mx276 
  // BSIM@ covered_modules=1 :   NAND3_X0P5A_A12TR c0nm_b0m_v0m_u80 (.A(c0nm_b0m_v0m_n95), .B(c0nm_b0m_v0m_n94), .C(c0nm_b0m_v0m_n72), .Y(c0nm_b0m_v0m_n100));
  // BSIM@ modules: mx167 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0nm_b0m_v0m_u68 (.A0(c0nm_b0m_v0m_n99), .A1(c0nm_b0m_v0m_n31), .B0(c0nm_b0m_v0m_n100), .B1(c0nm_b0m_v0m_n32), .C0(reset), .Y(c0nm_b0m_v0m_n101));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR c0nm_b0m_v0m_u82 (.A(c0nm_b0m_v0m_n99), .B(c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n102));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u79 (.A(c0nm_b0m_v0m_n98), .B(c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_n100), .Y(c0nm_b0m_v0m_n103));
  // BSIM@ modules: mx309 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u176 (.A(c0nm_b0m_v0m_n192), .Y(c0nm_b0m_v0m_n104));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u275 (.A(c0nm_b0m_v0m_buffers2_0_), .Y(c0nm_b0m_v0m_n105));
  // BSIM@ modules: mx366 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0nm_b0m_v0m_u85 (.A0(c0nm_b0m_v0m_n108), .A1(c0nm_b0m_v0m_n25), .B0(c0nm_b0m_v0m_n109), .B1(c0nm_b0m_v0m_n27), .C0(reset), .Y(c0nm_b0m_v0m_n106));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u167 (.A(c0nm_b0m_v0m_n187), .B(c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_n94), .Y(c0nm_b0m_v0m_n107));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u179 (.A(c0nm_b0m_v0m_n94), .Y(c0nm_b0m_v0m_n108));
  // BSIM@ modules: mx276 
  // BSIM@ covered_modules=1 :   NAND3_X0P5A_A12TR c0nm_b0m_v0m_u164 (.A(c0nm_b0m_v0m_n93), .B(c0nm_b0m_v0m_n95), .C(c0nm_b0m_v0m_n72), .Y(c0nm_b0m_v0m_n109));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0nm_b0m_v0m_u209 (.A(debitout_0), .B(reset), .Y(c0nm_b0m_v0m_n11));
  // BSIM@ modules: mx309 
  // BSIM@ covered_modules=1 :   OR2_X0P5M_A12TR c0nm_b0m_v0m_u173 (.A(c0nm_b0m_v0m_n187), .B(debitout_0), .Y(c0nm_b0m_v0m_n110));
  NAND4_X0P5A_A12TR c0nm_b0m_v0m_u174 (.A(c0nm_b0m_v0m_n96), .B(c0nm_b0m_v0m_n104), .C(c0nm_b0m_v0m_n187), .D(c0nm_v0m_n9), .Y(c0nm_b0m_v0m_n111));
  // BSIM@ modules: mx400 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0nm_b0m_v0m_u87 (.A0(c0nm_b0m_v0m_n113), .A1(c0nm_b0m_v0m_n114), .B0(c0nm_b0m_v0m_buffers0_0_), .B1(c0nm_b0m_v0m_n115), .C0(debitout_0), .Y(c0nm_b0m_v0m_n112));
  // BSIM@ modules: mx309 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0nm_b0m_v0m_u171 (.A(c0nm_b0m_v0m_n104), .B(debitout_0), .Y(c0nm_b0m_v0m_n113));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u270 (.A(c0nm_b0m_v0m_n61), .Y(c0nm_b0m_v0m_n114));
  // BSIM@ modules: mx309 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0nm_b0m_v0m_u172 (.A(c0nm_b0m_v0m_n96), .B(debitout_0), .Y(c0nm_b0m_v0m_n115));
  // BSIM@ modules: mx336 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u98 (.A(c0nm_b0m_v0m_n128), .Y(c0nm_b0m_v0m_n116));
  // BSIM@ modules: mx53 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u90 (.A0(c0nm_b0m_v0m_buffers0_0_), .A1(c0nm_b0m_v0m_n120), .B0(c0nm_b0m_v0m_buffers2_0_), .B1(c0nm_b0m_v0m_n121), .Y(c0nm_b0m_v0m_n117));
  // BSIM@ modules: mx30 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u89 (.A0(c0nm_b0m_v0m_n119), .A1(c0nm_b0m_v0m_n114), .B0(flitin_0[0]), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n118));
  // BSIM@ modules: mx336 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0nm_b0m_v0m_u191 (.A(c0nm_b0m_v0m_n93), .B(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n119));
  AOI21_X0P5M_A12TR c0nm_b0m_v0m_u16 (.A0(c0nm_b0m_v0m_n4), .A1(c0nm_b0m_v0m_n16), .B0(c0nm_b0m_v0m_n11), .Y(c0nm_b0m_v0m_n12));
  // BSIM@ modules: mx354 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0nm_b0m_v0m_u185 (.A(c0nm_b0m_v0m_n95), .B(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n120));
  // BSIM@ modules: mx354 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0nm_b0m_v0m_u187 (.A(c0nm_b0m_v0m_n94), .B(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n121));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u267 (.A(c0nm_b0m_v0m_buffers2_1_), .Y(c0nm_b0m_v0m_n122));
  // BSIM@ modules: mx366 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0nm_b0m_v0m_u92 (.A0(c0nm_b0m_v0m_n108), .A1(c0nm_b0m_v0m_n31), .B0(c0nm_b0m_v0m_n109), .B1(c0nm_b0m_v0m_n32), .C0(reset), .Y(c0nm_b0m_v0m_n123));
  // BSIM@ modules: mx401 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0nm_b0m_v0m_u94 (.A0(c0nm_b0m_v0m_n113), .A1(c0nm_b0m_v0m_n125), .B0(c0nm_b0m_v0m_buffers0_1_), .B1(c0nm_b0m_v0m_n115), .C0(debitout_0), .Y(c0nm_b0m_v0m_n124));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u265 (.A(c0nm_b0m_v0m_n60), .Y(c0nm_b0m_v0m_n125));
  // BSIM@ modules: mx53 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u97 (.A0(c0nm_b0m_v0m_buffers0_1_), .A1(c0nm_b0m_v0m_n120), .B0(c0nm_b0m_v0m_buffers2_1_), .B1(c0nm_b0m_v0m_n121), .Y(c0nm_b0m_v0m_n126));
  // BSIM@ modules: mx30 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u96 (.A0(c0nm_b0m_v0m_n119), .A1(c0nm_b0m_v0m_n125), .B0(flitin_0[1]), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n127));
  // BSIM@ modules: mx336 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0nm_b0m_v0m_u182 (.A(c0nm_b0m_v0m_n28), .B(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n128));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR c0nm_b0m_v0m_u178 (.A(c0nm_b0m_v0m_n108), .B(c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n129));
  NAND2_X0P5A_A12TR c0nm_b0m_v0m_u14 (.A(c0nm_b0m_v0m_n10), .B(c0nm_b0m_v0m_head_0_), .Y(c0nm_b0m_v0m_n13));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u163 (.A(c0nm_b0m_v0m_n107), .B(c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_n109), .Y(c0nm_b0m_v0m_n130));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u249 (.A(c0nm_b0m_v0m_buffers2_2_), .Y(c0nm_b0m_v0m_n131));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u101 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n35), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n131), .C0(c0nm_b0m_v0m_n133), .Y(c0nm_b0m_v0m_n132));
  // BSIM@ modules: mx64 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u102 (.A0(c0nm_b0m_v0m_buffers0_2_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n134), .Y(c0nm_b0m_v0m_n133));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u247 (.A(c0nm_b0m_v0m_n59), .Y(c0nm_b0m_v0m_n134));
  // BSIM@ modules: mx336 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u190 (.A(c0nm_b0m_v0m_n119), .Y(c0nm_b0m_v0m_n135));
  // BSIM@ modules: mx53 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u105 (.A0(c0nm_b0m_v0m_buffers2_2_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_2_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n136));
  // BSIM@ modules: mx31 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u104 (.A0(c0nm_b0m_v0m_buffers3_2_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_2_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n137));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u244 (.A(c0nm_b0m_v0m_buffers2_3_), .Y(c0nm_b0m_v0m_n138));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u108 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n38), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n138), .C0(c0nm_b0m_v0m_n140), .Y(c0nm_b0m_v0m_n139));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u13 (.A(c0nm_b0m_v0m_head_1_), .Y(c0nm_b0m_v0m_n14));
  // BSIM@ modules: mx64 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u109 (.A0(c0nm_b0m_v0m_buffers0_3_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n141), .Y(c0nm_b0m_v0m_n140));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u242 (.A(c0nm_b0m_v0m_n58), .Y(c0nm_b0m_v0m_n141));
  // BSIM@ modules: mx53 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u112 (.A0(c0nm_b0m_v0m_buffers2_3_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_3_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n142));
  // BSIM@ modules: mx31 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u111 (.A0(c0nm_b0m_v0m_buffers3_3_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_3_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n143));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u239 (.A(c0nm_b0m_v0m_buffers2_4_), .Y(c0nm_b0m_v0m_n144));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u115 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n41), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n144), .C0(c0nm_b0m_v0m_n146), .Y(c0nm_b0m_v0m_n145));
  // BSIM@ modules: mx64 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u116 (.A0(c0nm_b0m_v0m_buffers0_4_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n147), .Y(c0nm_b0m_v0m_n146));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u237 (.A(c0nm_b0m_v0m_n57), .Y(c0nm_b0m_v0m_n147));
  // BSIM@ modules: mx53 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u119 (.A0(c0nm_b0m_v0m_buffers2_4_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_4_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n148));
  // BSIM@ modules: mx31 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u118 (.A0(c0nm_b0m_v0m_buffers3_4_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_4_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n149));
  // BSIM@ modules: mx309 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u277 (.A(c0nm_b0m_v0m_head_2_), .Y(c0nm_b0m_v0m_n15));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u234 (.A(c0nm_b0m_v0m_buffers2_5_), .Y(c0nm_b0m_v0m_n150));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u122 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n44), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n150), .C0(c0nm_b0m_v0m_n152), .Y(c0nm_b0m_v0m_n151));
  // BSIM@ modules: mx64 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u123 (.A0(c0nm_b0m_v0m_buffers0_5_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n153), .Y(c0nm_b0m_v0m_n152));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u232 (.A(c0nm_b0m_v0m_n56), .Y(c0nm_b0m_v0m_n153));
  // BSIM@ modules: mx53 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u126 (.A0(c0nm_b0m_v0m_buffers2_5_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_5_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n154));
  // BSIM@ modules: mx31 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u125 (.A0(c0nm_b0m_v0m_buffers3_5_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_5_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n155));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u229 (.A(c0nm_b0m_v0m_buffers2_6_), .Y(c0nm_b0m_v0m_n156));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u129 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n47), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n156), .C0(c0nm_b0m_v0m_n158), .Y(c0nm_b0m_v0m_n157));
  // BSIM@ modules: mx64 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u130 (.A0(c0nm_b0m_v0m_buffers0_6_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n159), .Y(c0nm_b0m_v0m_n158));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u227 (.A(c0nm_b0m_v0m_n55), .Y(c0nm_b0m_v0m_n159));
  // BSIM@ modules: mx309 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u278 (.A(c0nm_b0m_v0m_head_0_), .Y(c0nm_b0m_v0m_n16));
  // BSIM@ modules: mx53 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u133 (.A0(c0nm_b0m_v0m_buffers2_6_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_6_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n160));
  // BSIM@ modules: mx31 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u132 (.A0(c0nm_b0m_v0m_buffers3_6_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_6_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n161));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u224 (.A(c0nm_b0m_v0m_buffers2_7_), .Y(c0nm_b0m_v0m_n162));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u136 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n62), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n162), .C0(c0nm_b0m_v0m_n164), .Y(c0nm_b0m_v0m_n163));
  // BSIM@ modules: mx64 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u137 (.A0(c0nm_b0m_v0m_buffers0_7_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n165), .Y(c0nm_b0m_v0m_n164));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u222 (.A(c0nm_b0m_v0m_n54), .Y(c0nm_b0m_v0m_n165));
  // BSIM@ modules: mx53 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u140 (.A0(c0nm_b0m_v0m_buffers2_7_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_7_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n166));
  // BSIM@ modules: mx31 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u139 (.A0(c0nm_b0m_v0m_buffers3_7_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_7_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n167));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u219 (.A(c0nm_b0m_v0m_buffers2_8_), .Y(c0nm_b0m_v0m_n168));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u143 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n65), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n168), .C0(c0nm_b0m_v0m_n170), .Y(c0nm_b0m_v0m_n169));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u168 (.A(c0nm_b0m_v0m_n188), .Y(c0nm_b0m_v0m_n17));
  // BSIM@ modules: mx64 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u144 (.A0(c0nm_b0m_v0m_buffers0_8_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n171), .Y(c0nm_b0m_v0m_n170));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u217 (.A(c0nm_b0m_v0m_n53), .Y(c0nm_b0m_v0m_n171));
  AND4_X0P5M_A12TR c0nm_b0m_v0m_u260 (.A(debitout_0), .B(c0nm_headflit[0]), .C(c0nm_b0m_v0m_n264), .D(c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n1710));
  // BSIM@ modules: mx53 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u147 (.A0(c0nm_b0m_v0m_buffers2_8_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_8_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n172));
  // BSIM@ modules: mx31 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u146 (.A0(c0nm_b0m_v0m_buffers3_8_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_8_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n173));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u214 (.A(c0nm_b0m_v0m_buffers2_9_), .Y(c0nm_b0m_v0m_n174));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u150 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n68), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n174), .C0(c0nm_b0m_v0m_n176), .Y(c0nm_b0m_v0m_n175));
  // BSIM@ modules: mx64 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u151 (.A0(c0nm_b0m_v0m_buffers0_9_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n177), .Y(c0nm_b0m_v0m_n176));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u212 (.A(c0nm_b0m_v0m_n52), .Y(c0nm_b0m_v0m_n177));
  // BSIM@ modules: mx53 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u154 (.A0(c0nm_b0m_v0m_buffers2_9_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_9_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n178));
  // BSIM@ modules: mx31 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u153 (.A0(c0nm_b0m_v0m_buffers3_9_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_9_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n179));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u32 (.A(c0nm_b0m_v0m_n22), .B(c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_n28), .Y(c0nm_b0m_v0m_n18));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u259 (.A(c0nm_b0m_v0m_buffers2_10_), .Y(c0nm_b0m_v0m_n180));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u157 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n71), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n180), .C0(c0nm_b0m_v0m_n182), .Y(c0nm_b0m_v0m_n181));
  // BSIM@ modules: mx64 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u158 (.A0(c0nm_b0m_v0m_buffers0_10_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n183), .Y(c0nm_b0m_v0m_n182));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u257 (.A(c0nm_b0m_v0m_n51), .Y(c0nm_b0m_v0m_n183));
  // BSIM@ modules: mx53 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u161 (.A0(c0nm_b0m_v0m_buffers2_10_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_10_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n184));
  // BSIM@ modules: mx31 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u160 (.A0(c0nm_b0m_v0m_buffers3_10_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_10_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n185));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u254 (.A(c0nm_b0m_v0m_buffers2_11_), .Y(c0nm_b0m_v0m_n186));
  // BSIM@ modules: mx309 
  // BSIM@ covered_modules=1 :   NAND3_X0P5A_A12TR c0nm_b0m_v0m_u276 (.A(c0nm_b0m_v0m_n16), .B(c0nm_b0m_v0m_n15), .C(c0nm_b0m_v0m_head_1_), .Y(c0nm_b0m_v0m_n187));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u169 (.A0(c0nm_b0m_v0m_n21), .A1(c0nm_b0m_v0m_n111), .B0(c0nm_b0m_v0m_n186), .B1(c0nm_b0m_v0m_n110), .C0(c0nm_b0m_v0m_n189), .Y(c0nm_b0m_v0m_n188));
  // BSIM@ modules: mx64 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u170 (.A0(c0nm_b0m_v0m_n115), .A1(c0nm_b0m_v0m_buffers0_11_), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n190), .Y(c0nm_b0m_v0m_n189));
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u180 (.A0(c0nm_b0m_v0m_n50), .A1(c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n194), .C0(c0nm_b0m_v0m_n195), .Y(c0nm_b0m_v0m_n19));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u252 (.A(c0nm_b0m_v0m_n50), .Y(c0nm_b0m_v0m_n190));
  // BSIM@ modules: mx309 
  // BSIM@ covered_modules=1 :   NOR3_X0P5A_A12TR c0nm_b0m_v0m_u271 (.A(c0nm_b0m_v0m_head_1_), .B(c0nm_b0m_v0m_head_2_), .C(c0nm_b0m_v0m_n16), .Y(c0nm_b0m_v0m_n192));
  // BSIM@ modules: mx309 
  // BSIM@ covered_modules=1 :   NOR3_X0P5A_A12TR c0nm_b0m_v0m_u272 (.A(c0nm_b0m_v0m_head_1_), .B(c0nm_b0m_v0m_head_2_), .C(c0nm_b0m_v0m_head_0_), .Y(c0nm_b0m_v0m_n193));
  // BSIM@ modules: mx53 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u184 (.A0(c0nm_b0m_v0m_buffers2_11_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_11_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n194));
  // BSIM@ modules: mx31 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u181 (.A0(c0nm_b0m_v0m_buffers3_11_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_n1), .B1(c0nm_b0m_wdata_11_), .Y(c0nm_b0m_v0m_n195));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0nm_b0m_v0m_u207 (.A0(c0nm_b0m_rdata[11]), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_b0m_headflit_11_), .Y(c0nm_b0m_v0m_n196));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0nm_b0m_v0m_u206 (.A0(c0nm_b0m_rdata[10]), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_b0m_headflit_10_), .Y(c0nm_b0m_v0m_n197));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0nm_b0m_v0m_u205 (.A0(c0nm_b0m_rdata[9]), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_b0m_headflit_9_), .Y(c0nm_b0m_v0m_n198));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0nm_b0m_v0m_u204 (.A0(c0nm_b0m_rdata[8]), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_b0m_headflit_8_), .Y(c0nm_b0m_v0m_n199));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR c0nm_b0m_v0m_u4 (.A(c0nm_b0m_v0m_n1), .B(c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n2));
  // BSIM@ modules: mx346 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR c0nm_b0m_v0m_u31 (.A(c0nm_b0m_v0m_n26), .B(c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n20));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0nm_b0m_v0m_u203 (.A0(c0nm_b0m_rdata[7]), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit[7]), .Y(c0nm_b0m_v0m_n200));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0nm_b0m_v0m_u202 (.A0(c0nm_b0m_rdata[6]), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit[6]), .Y(c0nm_b0m_v0m_n201));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0nm_b0m_v0m_u201 (.A0(c0nm_b0m_rdata[5]), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit[5]), .Y(c0nm_b0m_v0m_n202));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0nm_b0m_v0m_u200 (.A0(c0nm_b0m_rdata[4]), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit[4]), .Y(c0nm_b0m_v0m_n203));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0nm_b0m_v0m_u199 (.A0(c0nm_b0m_rdata[3]), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit[3]), .Y(c0nm_b0m_v0m_n204));
  // BSIM@ modules: mx249 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0nm_b0m_v0m_u198 (.A0(c0nm_b0m_rdata[2]), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit[2]), .Y(c0nm_b0m_v0m_n205));
  // BSIM@ modules: mx245 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR c0nm_b0m_v0m_u196 (.A(c0nm_b0m_v0m_n263), .B(c0nm_b0m_rdata[1]), .S0(c0nm_b0m_v0m_n11), .Y(c0nm_b0m_v0m_n206));
  // BSIM@ modules: mx245 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR c0nm_b0m_v0m_u194 (.A(c0nm_b0m_v0m_n262), .B(c0nm_b0m_rdata[0]), .S0(c0nm_b0m_v0m_n11), .Y(c0nm_b0m_v0m_n207));
  // BSIM@ modules: mx102 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u162 (.A0(c0nm_b0m_v0m_n19), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n17), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n186), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n208));
  // BSIM@ modules: mx102 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u155 (.A0(c0nm_b0m_v0m_n70), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n69), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n180), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n209));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u253 (.A(c0nm_b0m_v0m_buffers3_11_), .Y(c0nm_b0m_v0m_n21));
  // BSIM@ modules: mx102 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u148 (.A0(c0nm_b0m_v0m_n67), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n66), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n174), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n210));
  // BSIM@ modules: mx102 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u141 (.A0(c0nm_b0m_v0m_n64), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n63), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n168), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n211));
  // BSIM@ modules: mx102 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u134 (.A0(c0nm_b0m_v0m_n49), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n48), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n162), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n212));
  // BSIM@ modules: mx102 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u127 (.A0(c0nm_b0m_v0m_n46), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n45), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n156), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n213));
  // BSIM@ modules: mx102 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u120 (.A0(c0nm_b0m_v0m_n43), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n42), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n150), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n214));
  // BSIM@ modules: mx102 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u113 (.A0(c0nm_b0m_v0m_n40), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n39), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n144), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n215));
  // BSIM@ modules: mx102 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u106 (.A0(c0nm_b0m_v0m_n37), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n36), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n138), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n216));
  // BSIM@ modules: mx102 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u99 (.A0(c0nm_b0m_v0m_n34), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n33), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n131), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n217));
  // BSIM@ modules: mx366 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u91 (.A(c0nm_b0m_v0m_n122), .B(c0nm_b0m_v0m_n123), .S0(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n218));
  // BSIM@ modules: mx366 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u84 (.A(c0nm_b0m_v0m_n105), .B(c0nm_b0m_v0m_n106), .S0(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n219));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u33 (.A(c0nm_b0m_v0m_n72), .B(c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_n73), .Y(c0nm_b0m_v0m_n22));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u78 (.A0(c0nm_b0m_v0m_n19), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n17), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n50), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n220));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u77 (.A0(c0nm_b0m_v0m_n70), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n69), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n51), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n221));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u76 (.A0(c0nm_b0m_v0m_n67), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n66), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n52), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n222));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u75 (.A0(c0nm_b0m_v0m_n64), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n63), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n53), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n223));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u74 (.A0(c0nm_b0m_v0m_n49), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n48), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n54), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n224));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u73 (.A0(c0nm_b0m_v0m_n46), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n45), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n55), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n225));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u72 (.A0(c0nm_b0m_v0m_n43), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n42), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n56), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n226));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u71 (.A0(c0nm_b0m_v0m_n40), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n39), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n57), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n227));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u70 (.A0(c0nm_b0m_v0m_n37), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n36), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n58), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n228));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u69 (.A0(c0nm_b0m_v0m_n34), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n33), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n59), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n229));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u273 (.A(c0nm_b0m_v0m_buffers3_0_), .Y(c0nm_b0m_v0m_n23));
  // BSIM@ modules: mx247 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u67 (.A(c0nm_b0m_v0m_n60), .B(c0nm_b0m_v0m_n101), .S0(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n230));
  // BSIM@ modules: mx247 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u65 (.A(c0nm_b0m_v0m_n61), .B(c0nm_b0m_v0m_n97), .S0(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n231));
  // BSIM@ modules: mx104 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u58 (.A0(c0nm_b0m_v0m_n19), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n17), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n92), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n232));
  // BSIM@ modules: mx104 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u56 (.A0(c0nm_b0m_v0m_n70), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n69), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n91), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n233));
  // BSIM@ modules: mx104 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u54 (.A0(c0nm_b0m_v0m_n67), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n66), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n90), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n234));
  // BSIM@ modules: mx104 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u52 (.A0(c0nm_b0m_v0m_n64), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n63), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n89), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n235));
  // BSIM@ modules: mx104 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u50 (.A0(c0nm_b0m_v0m_n49), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n48), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n88), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n236));
  // BSIM@ modules: mx104 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u48 (.A0(c0nm_b0m_v0m_n46), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n45), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n87), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n237));
  // BSIM@ modules: mx104 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u46 (.A0(c0nm_b0m_v0m_n43), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n42), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n86), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n238));
  // BSIM@ modules: mx104 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u44 (.A0(c0nm_b0m_v0m_n40), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n39), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n85), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n239));
  // BSIM@ modules: mx369 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0nm_b0m_v0m_u19 (.A0(c0nm_b0m_v0m_n25), .A1(c0nm_b0m_v0m_n26), .B0(c0nm_b0m_v0m_n27), .B1(c0nm_b0m_v0m_n28), .C0(reset), .Y(c0nm_b0m_v0m_n24));
  // BSIM@ modules: mx104 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u42 (.A0(c0nm_b0m_v0m_n37), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n36), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n84), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n240));
  // BSIM@ modules: mx104 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u40 (.A0(c0nm_b0m_v0m_n34), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n33), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n83), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n241));
  // BSIM@ modules: mx368 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u37 (.A(c0nm_b0m_v0m_n79), .B(c0nm_b0m_v0m_n80), .S0(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n242));
  // BSIM@ modules: mx368 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u34 (.A(c0nm_b0m_v0m_n74), .B(c0nm_b0m_v0m_n75), .S0(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n243));
  // BSIM@ modules: mx105 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u30 (.A0(c0nm_b0m_v0m_n69), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n70), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n71), .Y(c0nm_b0m_v0m_n244));
  // BSIM@ modules: mx105 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u29 (.A0(c0nm_b0m_v0m_n66), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n67), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n68), .Y(c0nm_b0m_v0m_n245));
  // BSIM@ modules: mx105 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u28 (.A0(c0nm_b0m_v0m_n63), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n64), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n65), .Y(c0nm_b0m_v0m_n246));
  // BSIM@ modules: mx105 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u27 (.A0(c0nm_b0m_v0m_n48), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n49), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n62), .Y(c0nm_b0m_v0m_n247));
  // BSIM@ modules: mx105 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u26 (.A0(c0nm_b0m_v0m_n45), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n46), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n47), .Y(c0nm_b0m_v0m_n248));
  // BSIM@ modules: mx105 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u25 (.A0(c0nm_b0m_v0m_n42), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n43), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n44), .Y(c0nm_b0m_v0m_n249));
  OAI211_X0P5M_A12TR c0nm_b0m_v0m_u88 (.A0(c0nm_b0m_v0m_n116), .A1(c0nm_b0m_v0m_n23), .B0(c0nm_b0m_v0m_n117), .C0(c0nm_b0m_v0m_n118), .Y(c0nm_b0m_v0m_n25));
  // BSIM@ modules: mx105 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u24 (.A0(c0nm_b0m_v0m_n39), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n40), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n41), .Y(c0nm_b0m_v0m_n250));
  // BSIM@ modules: mx105 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u23 (.A0(c0nm_b0m_v0m_n36), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n37), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n38), .Y(c0nm_b0m_v0m_n251));
  // BSIM@ modules: mx105 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u22 (.A0(c0nm_b0m_v0m_n33), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n34), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n35), .Y(c0nm_b0m_v0m_n252));
  // BSIM@ modules: mx369 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u20 (.A(c0nm_b0m_v0m_n29), .B(c0nm_b0m_v0m_n30), .S0(c0nm_b0m_v0m_n22), .Y(c0nm_b0m_v0m_n253));
  // BSIM@ modules: mx369 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u18 (.A(c0nm_b0m_v0m_n23), .B(c0nm_b0m_v0m_n24), .S0(c0nm_b0m_v0m_n22), .Y(c0nm_b0m_v0m_n254));
  // BSIM@ modules: mx105 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0nm_b0m_v0m_u17 (.A0(c0nm_b0m_v0m_n17), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n19), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n21), .C1(c0nm_b0m_v0m_n22), .Y(c0nm_b0m_v0m_n255));
  OA21A1OI2_X0P5M_A12TR c0nm_b0m_v0m_u15 (.A0(reset), .A1(c0nm_b0m_v0m_head_1_), .B0(c0nm_b0m_v0m_n12), .C0(c0nm_b0m_v0m_n15), .Y(c0nm_b0m_v0m_n256));
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u12 (.A(c0nm_b0m_v0m_n12), .B(c0nm_b0m_v0m_n13), .S0(c0nm_b0m_v0m_n14), .Y(c0nm_b0m_v0m_n257));
  MXT2_X0P5M_A12TR c0nm_b0m_v0m_u11 (.A(c0nm_b0m_v0m_n10), .B(c0nm_b0m_v0m_n11), .S0(c0nm_b0m_v0m_head_0_), .Y(c0nm_b0m_v0m_n258));
  OA21A1OI2_X0P5M_A12TR c0nm_b0m_v0m_u8 (.A0(c0nm_b0m_v0m_tail_1_), .A1(reset), .B0(c0nm_b0m_v0m_n5), .C0(c0nm_b0m_v0m_n9), .Y(c0nm_b0m_v0m_n259));
  // BSIM@ modules: mx276 
  // BSIM@ covered_modules=1 :   OAI21_X0P5M_A12TR c0nm_b0m_v0m_u166 (.A0(c0nm_b0m_v0m_n3), .A1(c0nm_b0m_v0m_n7), .B0(c0nm_b0m_v0m_n9), .Y(c0nm_b0m_v0m_n26));
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u5 (.A(c0nm_b0m_v0m_n5), .B(c0nm_b0m_v0m_n6), .S0(c0nm_b0m_v0m_n7), .Y(c0nm_b0m_v0m_n260));
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u3 (.A(c0nm_b0m_v0m_n1), .B(c0nm_b0m_v0m_n2), .S0(c0nm_b0m_v0m_n3), .Y(c0nm_b0m_v0m_n261));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   NAND2B_X0P5M_A12TR c0nm_b0m_v0m_u195 (.AN(c0nm_headflit[0]), .B(c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n262));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR c0nm_b0m_v0m_u197 (.A(c0nm_b0m_v0m_n264), .B(c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n263));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u262 (.A(c0nm_headflit[1]), .Y(c0nm_b0m_v0m_n264));
  // BSIM@ modules: mx374 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u211 (.A0(c0nm_b0m_v0m_buffers0_9_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n177), .Y(c0nm_b0m_v0m_n265));
  // BSIM@ modules: mx374 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u216 (.A0(c0nm_b0m_v0m_buffers0_8_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n171), .Y(c0nm_b0m_v0m_n266));
  // BSIM@ modules: mx374 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u221 (.A0(c0nm_b0m_v0m_buffers0_7_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n165), .Y(c0nm_b0m_v0m_n267));
  // BSIM@ modules: mx42 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u226 (.A0(c0nm_b0m_v0m_buffers0_6_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n159), .Y(c0nm_b0m_v0m_n268));
  // BSIM@ modules: mx42 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u231 (.A0(c0nm_b0m_v0m_buffers0_5_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n153), .Y(c0nm_b0m_v0m_n269));
  // BSIM@ modules: mx400 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u86 (.A0(c0nm_b0m_v0m_n110), .A1(c0nm_b0m_v0m_n105), .B0(c0nm_b0m_v0m_n111), .B1(c0nm_b0m_v0m_n23), .C0(c0nm_b0m_v0m_n112), .Y(c0nm_b0m_v0m_n27));
  // BSIM@ modules: mx374 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u236 (.A0(c0nm_b0m_v0m_buffers0_4_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n147), .Y(c0nm_b0m_v0m_n270));
  // BSIM@ modules: mx42 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u241 (.A0(c0nm_b0m_v0m_buffers0_3_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n141), .Y(c0nm_b0m_v0m_n271));
  // BSIM@ modules: mx374 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u246 (.A0(c0nm_b0m_v0m_buffers0_2_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n134), .Y(c0nm_b0m_v0m_n272));
  // BSIM@ modules: mx374 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u251 (.A0(c0nm_b0m_v0m_n193), .A1(c0nm_b0m_v0m_buffers0_11_), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n190), .Y(c0nm_b0m_v0m_n273));
  // BSIM@ modules: mx374 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u256 (.A0(c0nm_b0m_v0m_buffers0_10_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n183), .Y(c0nm_b0m_v0m_n274));
  // BSIM@ modules: mx42 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u264 (.A0(c0nm_b0m_v0m_buffers0_1_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n125), .Y(c0nm_b0m_v0m_n275));
  // BSIM@ modules: mx42 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_b0m_v0m_u269 (.A0(c0nm_b0m_v0m_buffers0_0_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n114), .Y(c0nm_b0m_v0m_n276));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u183 (.A(c0nm_b0m_v0m_n95), .B(c0nm_b0m_v0m_n94), .C(c0nm_b0m_v0m_n93), .Y(c0nm_b0m_v0m_n28));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u266 (.A(c0nm_b0m_v0m_buffers3_1_), .Y(c0nm_b0m_v0m_n29));
  // BSIM@ modules: mx276 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u189 (.A(c0nm_b0m_v0m_tail_0_), .Y(c0nm_b0m_v0m_n3));
  // BSIM@ modules: mx369 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0nm_b0m_v0m_u21 (.A0(c0nm_b0m_v0m_n31), .A1(c0nm_b0m_v0m_n26), .B0(c0nm_b0m_v0m_n32), .B1(c0nm_b0m_v0m_n28), .C0(reset), .Y(c0nm_b0m_v0m_n30));
  OAI211_X0P5M_A12TR c0nm_b0m_v0m_u95 (.A0(c0nm_b0m_v0m_n116), .A1(c0nm_b0m_v0m_n29), .B0(c0nm_b0m_v0m_n126), .C0(c0nm_b0m_v0m_n127), .Y(c0nm_b0m_v0m_n31));
  // BSIM@ modules: mx401 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u93 (.A0(c0nm_b0m_v0m_n110), .A1(c0nm_b0m_v0m_n122), .B0(c0nm_b0m_v0m_n111), .B1(c0nm_b0m_v0m_n29), .C0(c0nm_b0m_v0m_n124), .Y(c0nm_b0m_v0m_n32));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u100 (.A(c0nm_b0m_v0m_n132), .Y(c0nm_b0m_v0m_n33));
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u103 (.A0(c0nm_b0m_v0m_n59), .A1(c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n136), .C0(c0nm_b0m_v0m_n137), .Y(c0nm_b0m_v0m_n34));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u248 (.A(c0nm_b0m_v0m_buffers3_2_), .Y(c0nm_b0m_v0m_n35));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u107 (.A(c0nm_b0m_v0m_n139), .Y(c0nm_b0m_v0m_n36));
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u110 (.A0(c0nm_b0m_v0m_n58), .A1(c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n142), .C0(c0nm_b0m_v0m_n143), .Y(c0nm_b0m_v0m_n37));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u243 (.A(c0nm_b0m_v0m_buffers3_3_), .Y(c0nm_b0m_v0m_n38));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u114 (.A(c0nm_b0m_v0m_n145), .Y(c0nm_b0m_v0m_n39));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u261 (.A(reset), .Y(c0nm_b0m_v0m_n4));
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u117 (.A0(c0nm_b0m_v0m_n57), .A1(c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n148), .C0(c0nm_b0m_v0m_n149), .Y(c0nm_b0m_v0m_n40));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u238 (.A(c0nm_b0m_v0m_buffers3_4_), .Y(c0nm_b0m_v0m_n41));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u121 (.A(c0nm_b0m_v0m_n151), .Y(c0nm_b0m_v0m_n42));
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u124 (.A0(c0nm_b0m_v0m_n56), .A1(c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n154), .C0(c0nm_b0m_v0m_n155), .Y(c0nm_b0m_v0m_n43));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u233 (.A(c0nm_b0m_v0m_buffers3_5_), .Y(c0nm_b0m_v0m_n44));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u128 (.A(c0nm_b0m_v0m_n157), .Y(c0nm_b0m_v0m_n45));
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u131 (.A0(c0nm_b0m_v0m_n55), .A1(c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n160), .C0(c0nm_b0m_v0m_n161), .Y(c0nm_b0m_v0m_n46));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u228 (.A(c0nm_b0m_v0m_buffers3_6_), .Y(c0nm_b0m_v0m_n47));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u135 (.A(c0nm_b0m_v0m_n163), .Y(c0nm_b0m_v0m_n48));
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u138 (.A0(c0nm_b0m_v0m_n54), .A1(c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n166), .C0(c0nm_b0m_v0m_n167), .Y(c0nm_b0m_v0m_n49));
  AOI21_X0P5M_A12TR c0nm_b0m_v0m_u9 (.A0(c0nm_b0m_v0m_n3), .A1(c0nm_b0m_v0m_n4), .B0(c0nm_b0m_v0m_n8), .Y(c0nm_b0m_v0m_n5));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_11_ (.CK(clk), .QN(c0nm_b0m_v0m_n50), .D(c0nm_b0m_v0m_n220));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_10_ (.CK(clk), .QN(c0nm_b0m_v0m_n51), .D(c0nm_b0m_v0m_n221));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_9_ (.CK(clk), .QN(c0nm_b0m_v0m_n52), .D(c0nm_b0m_v0m_n222));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_8_ (.CK(clk), .QN(c0nm_b0m_v0m_n53), .D(c0nm_b0m_v0m_n223));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_7_ (.CK(clk), .QN(c0nm_b0m_v0m_n54), .D(c0nm_b0m_v0m_n224));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_6_ (.CK(clk), .QN(c0nm_b0m_v0m_n55), .D(c0nm_b0m_v0m_n225));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_5_ (.CK(clk), .QN(c0nm_b0m_v0m_n56), .D(c0nm_b0m_v0m_n226));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_4_ (.CK(clk), .QN(c0nm_b0m_v0m_n57), .D(c0nm_b0m_v0m_n227));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_3_ (.CK(clk), .QN(c0nm_b0m_v0m_n58), .D(c0nm_b0m_v0m_n228));
  // BSIM@ modules: mx251 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_2_ (.CK(clk), .QN(c0nm_b0m_v0m_n59), .D(c0nm_b0m_v0m_n229));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u6 (.A(c0nm_b0m_v0m_n1), .B(c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_tail_0_), .Y(c0nm_b0m_v0m_n6));
  // BSIM@ modules: mx247 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_1_ (.CK(clk), .QN(c0nm_b0m_v0m_n60), .D(c0nm_b0m_v0m_n230));
  // BSIM@ modules: mx247 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_0_ (.CK(clk), .QN(c0nm_b0m_v0m_n61), .D(c0nm_b0m_v0m_n231));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u223 (.A(c0nm_b0m_v0m_buffers3_7_), .Y(c0nm_b0m_v0m_n62));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u142 (.A(c0nm_b0m_v0m_n169), .Y(c0nm_b0m_v0m_n63));
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u145 (.A0(c0nm_b0m_v0m_n53), .A1(c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n172), .C0(c0nm_b0m_v0m_n173), .Y(c0nm_b0m_v0m_n64));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u218 (.A(c0nm_b0m_v0m_buffers3_8_), .Y(c0nm_b0m_v0m_n65));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u149 (.A(c0nm_b0m_v0m_n175), .Y(c0nm_b0m_v0m_n66));
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u152 (.A0(c0nm_b0m_v0m_n52), .A1(c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n178), .C0(c0nm_b0m_v0m_n179), .Y(c0nm_b0m_v0m_n67));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u213 (.A(c0nm_b0m_v0m_buffers3_9_), .Y(c0nm_b0m_v0m_n68));
  // BSIM@ modules: mx211 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u156 (.A(c0nm_b0m_v0m_n181), .Y(c0nm_b0m_v0m_n69));
  // BSIM@ modules: mx276 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u193 (.A(c0nm_b0m_v0m_tail_1_), .Y(c0nm_b0m_v0m_n7));
  OA211_X0P5M_A12TR c0nm_b0m_v0m_u159 (.A0(c0nm_b0m_v0m_n51), .A1(c0nm_b0m_v0m_n135), .B0(c0nm_b0m_v0m_n184), .C0(c0nm_b0m_v0m_n185), .Y(c0nm_b0m_v0m_n70));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u258 (.A(c0nm_b0m_v0m_buffers3_10_), .Y(c0nm_b0m_v0m_n71));
  // BSIM@ modules: mx276 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u165 (.A(c0nm_b0m_v0m_n26), .Y(c0nm_b0m_v0m_n72));
  AOI21_X0P5M_A12TR c0nm_b0m_v0m_u274 (.A0(c0nm_b0m_v0m_head_0_), .A1(c0nm_b0m_v0m_head_1_), .B0(c0nm_b0m_v0m_head_2_), .Y(c0nm_b0m_v0m_n73));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u36 (.A(c0nm_b0m_v0m_buffers0_0_), .Y(c0nm_b0m_v0m_n74));
  // BSIM@ modules: mx368 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0nm_b0m_v0m_u35 (.A0(c0nm_b0m_v0m_n77), .A1(c0nm_b0m_v0m_n25), .B0(c0nm_b0m_v0m_n78), .B1(c0nm_b0m_v0m_n27), .C0(reset), .Y(c0nm_b0m_v0m_n75));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u62 (.A(c0nm_b0m_v0m_n95), .B(c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_n96), .Y(c0nm_b0m_v0m_n76));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u64 (.A(c0nm_b0m_v0m_n95), .Y(c0nm_b0m_v0m_n77));
  // BSIM@ modules: mx276 
  // BSIM@ covered_modules=1 :   NAND3_X0P5A_A12TR c0nm_b0m_v0m_u61 (.A(c0nm_b0m_v0m_n93), .B(c0nm_b0m_v0m_n94), .C(c0nm_b0m_v0m_n72), .Y(c0nm_b0m_v0m_n78));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u39 (.A(c0nm_b0m_v0m_buffers0_1_), .Y(c0nm_b0m_v0m_n79));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0nm_b0m_v0m_u10 (.A(reset), .B(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n8));
  // BSIM@ modules: mx368 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0nm_b0m_v0m_u38 (.A0(c0nm_b0m_v0m_n77), .A1(c0nm_b0m_v0m_n31), .B0(c0nm_b0m_v0m_n78), .B1(c0nm_b0m_v0m_n32), .C0(reset), .Y(c0nm_b0m_v0m_n80));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR c0nm_b0m_v0m_u63 (.A(c0nm_b0m_v0m_n77), .B(c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n81));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u60 (.A(c0nm_b0m_v0m_n76), .B(c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_n78), .Y(c0nm_b0m_v0m_n82));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u41 (.A(c0nm_b0m_v0m_buffers0_2_), .Y(c0nm_b0m_v0m_n83));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u43 (.A(c0nm_b0m_v0m_buffers0_3_), .Y(c0nm_b0m_v0m_n84));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u45 (.A(c0nm_b0m_v0m_buffers0_4_), .Y(c0nm_b0m_v0m_n85));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u47 (.A(c0nm_b0m_v0m_buffers0_5_), .Y(c0nm_b0m_v0m_n86));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u49 (.A(c0nm_b0m_v0m_buffers0_6_), .Y(c0nm_b0m_v0m_n87));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u51 (.A(c0nm_b0m_v0m_buffers0_7_), .Y(c0nm_b0m_v0m_n88));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u53 (.A(c0nm_b0m_v0m_buffers0_8_), .Y(c0nm_b0m_v0m_n89));
  DFFQN_X1M_A12TR c0nm_b0m_v0m_tail_reg_2_ (.CK(clk), .QN(c0nm_b0m_v0m_n9), .D(c0nm_b0m_v0m_n259));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u55 (.A(c0nm_b0m_v0m_buffers0_9_), .Y(c0nm_b0m_v0m_n90));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u57 (.A(c0nm_b0m_v0m_buffers0_10_), .Y(c0nm_b0m_v0m_n91));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u59 (.A(c0nm_b0m_v0m_buffers0_11_), .Y(c0nm_b0m_v0m_n92));
  // BSIM@ modules: mx276 
  // BSIM@ covered_modules=1 :   NAND3_X0P5A_A12TR c0nm_b0m_v0m_u192 (.A(c0nm_b0m_v0m_tail_0_), .B(c0nm_b0m_v0m_n7), .C(c0nm_b0m_v0m_n9), .Y(c0nm_b0m_v0m_n93));
  // BSIM@ modules: mx276 
  // BSIM@ covered_modules=1 :   NAND3_X0P5A_A12TR c0nm_b0m_v0m_u188 (.A(c0nm_b0m_v0m_tail_1_), .B(c0nm_b0m_v0m_n3), .C(c0nm_b0m_v0m_n9), .Y(c0nm_b0m_v0m_n94));
  // BSIM@ modules: mx276 
  // BSIM@ covered_modules=1 :   NAND3_X0P5A_A12TR c0nm_b0m_v0m_u186 (.A(c0nm_b0m_v0m_n3), .B(c0nm_b0m_v0m_n7), .C(c0nm_b0m_v0m_n9), .Y(c0nm_b0m_v0m_n95));
  // BSIM@ modules: mx309 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u177 (.A(c0nm_b0m_v0m_n193), .Y(c0nm_b0m_v0m_n96));
  // BSIM@ modules: mx167 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0nm_b0m_v0m_u66 (.A0(c0nm_b0m_v0m_n99), .A1(c0nm_b0m_v0m_n25), .B0(c0nm_b0m_v0m_n100), .B1(c0nm_b0m_v0m_n27), .C0(reset), .Y(c0nm_b0m_v0m_n97));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u81 (.A(c0nm_b0m_v0m_n93), .B(c0nm_b0m_v0m_n4), .C(c0nm_b0m_v0m_n104), .Y(c0nm_b0m_v0m_n98));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_b0m_v0m_u83 (.A(c0nm_b0m_v0m_n93), .Y(c0nm_b0m_v0m_n99));
  // BSIM@ modules: mx405 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0nm_b0m_v0m_tail_reg_0_ (.CK(clk), .Q(c0nm_b0m_v0m_tail_0_), .D(c0nm_b0m_v0m_n261));
  // BSIM@ modules: mx405 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0nm_b0m_v0m_tail_reg_1_ (.CK(clk), .Q(c0nm_b0m_v0m_tail_1_), .D(c0nm_b0m_v0m_n260));
  // BSIM@ modules: mx320 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u13 (.A(flitin_0[10]), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_10_));
  // BSIM@ modules: mx320 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u12 (.A(flitin_0[11]), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_11_));
  // BSIM@ modules: mx320 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u11 (.A(flitin_0[2]), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_2_));
  // BSIM@ modules: mx320 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u10 (.A(flitin_0[3]), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_3_));
  // BSIM@ modules: mx320 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u9 (.A(flitin_0[4]), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_4_));
  // BSIM@ modules: mx320 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u8 (.A(flitin_0[5]), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_5_));
  // BSIM@ modules: mx320 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u7 (.A(flitin_0[6]), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_6_));
  // BSIM@ modules: mx320 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u6 (.A(flitin_0[7]), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_7_));
  // BSIM@ modules: mx320 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u5 (.A(flitin_0[8]), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_8_));
  // BSIM@ modules: mx320 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u4 (.A(flitin_0[9]), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_9_));
  // BSIM@ modules: mx400 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u268 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n105), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n23), .C0(c0nm_b0m_v0m_n276), .Y(c0nm_headflit[0]));
  // BSIM@ modules: mx401 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u263 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n122), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n29), .C0(c0nm_b0m_v0m_n275), .Y(c0nm_headflit[1]));
  // BSIM@ modules: mx374 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u245 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n131), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n35), .C0(c0nm_b0m_v0m_n272), .Y(c0nm_headflit[2]));
  // BSIM@ modules: mx207 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u240 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n138), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n38), .C0(c0nm_b0m_v0m_n271), .Y(c0nm_headflit[3]));
  // BSIM@ modules: mx374 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u235 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n144), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n41), .C0(c0nm_b0m_v0m_n270), .Y(c0nm_headflit[4]));
  // BSIM@ modules: mx207 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u230 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n150), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n44), .C0(c0nm_b0m_v0m_n269), .Y(c0nm_headflit[5]));
  // BSIM@ modules: mx207 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u225 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n156), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n47), .C0(c0nm_b0m_v0m_n268), .Y(c0nm_headflit[6]));
  // BSIM@ modules: mx374 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0nm_b0m_v0m_u220 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n162), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n62), .C0(c0nm_b0m_v0m_n267), .Y(c0nm_headflit[7]));
  NOR2B_X0P5M_A12TR c0nm_u4 (.AN(c0nm_headflit[1]), .B(c0nm_headflit[0]), .Y(c0nm_n1));
  // BSIM@ modules: mx343 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR c0nm_u3 (.A(flitin_0[1]), .B(flitin_0[0]), .Y(c0nm_n2));
  INV_X0P5B_A12TR c0nm_r0m_u6 (.A(c0nm_n1), .Y(c0nm_r0m_n1));
  AOI2XB1_X0P5M_A12TR c0nm_r0m_u10 (.A0(curry[2]), .A1N(c0nm_headflit[4]), .B0(c0nm_r0m_n11), .Y(c0nm_r0m_n10));
  NOR3_X0P5A_A12TR c0nm_r0m_u5 (.A(c0nm_r0m_n3), .B(reset), .C(c0nm_r0m_n1), .Y(c0nm_r0m_n100));
  AOI2XB1_X0P5M_A12TR c0nm_r0m_u11 (.A0(c0nm_headflit[4]), .A1N(curry[2]), .B0(c0nm_r0m_n12), .Y(c0nm_r0m_n11));
  NOR3_X0P5A_A12TR c0nm_r0m_u3 (.A(c0nm_r0m_n1), .B(reset), .C(c0nm_r0m_n2), .Y(c0nm_r0m_n110));
  // BSIM@ modules: mx29 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0nm_r0m_u12 (.A0(c0nm_r0m_n13), .A1(curry[0]), .B0(curry[1]), .B1(c0nm_r0m_n14), .Y(c0nm_r0m_n12));
  AOI2XB1_X0P5M_A12TR c0nm_r0m_u14 (.A0(c0nm_headflit[3]), .A1N(curry[1]), .B0(c0nm_headflit[2]), .Y(c0nm_r0m_n13));
  // BSIM@ modules: mx207 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_r0m_u13 (.A(c0nm_headflit[3]), .Y(c0nm_r0m_n14));
  // BSIM@ modules: mx334 
  // BSIM@ covered_modules=1 :   OR2_X0P5M_A12TR c0nm_r0m_u18 (.A(currx[0]), .B(c0nm_r0m_n9), .Y(c0nm_r0m_n15));
  // BSIM@ modules: mx319 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_r0m_u16 (.A(c0nm_r0m_n15), .B(currx[1]), .Y(c0nm_r0m_n16));
  INV_X0P5B_A12TR c0nm_r0m_u4 (.A(c0nm_r0m_n3), .Y(c0nm_r0m_n2));
  AO1B2_X0P5M_A12TR c0nm_r0m_u7 (.A0N(c0nm_r0m_n5), .B0(c0nm_r0m_n4), .B1(c0nm_headflit[7]), .Y(c0nm_r0m_n3));
  INV_X0P5B_A12TR c0nm_r0m_u20 (.A(currx[2]), .Y(c0nm_r0m_n4));
  OAI22_X0P5M_A12TR c0nm_r0m_u8 (.A0(c0nm_r0m_n6), .A1(c0nm_r0m_n7), .B0(c0nm_headflit[7]), .B1(c0nm_r0m_n4), .Y(c0nm_r0m_n5));
  OA21A1OI2_X0P5M_A12TR c0nm_r0m_u15 (.A0(currx[1]), .A1(c0nm_r0m_n15), .B0(c0nm_r0m_n8), .C0(c0nm_r0m_n16), .Y(c0nm_r0m_n6));
  // BSIM@ modules: mx110 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0nm_r0m_u9 (.A0(currx[1]), .A1(c0nm_r0m_n8), .B0(currx[0]), .B1(c0nm_r0m_n9), .C0(c0nm_r0m_n10), .Y(c0nm_r0m_n7));
  // BSIM@ modules: mx207 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_r0m_u17 (.A(c0nm_headflit[6]), .Y(c0nm_r0m_n8));
  // BSIM@ modules: mx207 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_r0m_u19 (.A(c0nm_headflit[5]), .Y(c0nm_r0m_n9));
  DFFQ_X1M_A12TR c0nm_r0m_vc_req_reg_0_ (.CK(clk), .Q(c0nm_routewire[0]), .D(c0nm_r0m_n100));
  DFFQ_X1M_A12TR c0nm_r0m_vc_req_reg_1_ (.CK(clk), .Q(c0nm_routewire[1]), .D(c0nm_r0m_n110));
  DFFQ_X1M_A12TR c0nm_v0m_full_reg (.CK(clk), .Q(c0nm_v0m_full), .D(c0nm_v0m_n64));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_v0m_u9 (.A(c0nm_v0m_n8), .Y(c0nm_v0m_n1));
  AOI32_X0P5M_A12TR c0nm_v0m_u12 (.A0(c0nm_v0m_n11), .A1(c0nm_v0m_n9), .A2(c0nm_n2), .B0(c0nm_v0m_full), .B1(c0nm_v0m_n12), .Y(c0nm_v0m_n10));
  INV_X0P5B_A12TR c0nm_v0m_u14 (.A(c0nm_v0m_n14), .Y(c0nm_v0m_n11));
  INV_X0P5B_A12TR c0nm_v0m_u13 (.A(c0nm_v0m_n13), .Y(c0nm_v0m_n12));
  // BSIM@ modules: mx356 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0nm_v0m_u30 (.A(c0nm_v0m_n9), .B(c0nm_n2), .Y(c0nm_v0m_n13));
  NAND3_X0P5A_A12TR c0nm_v0m_u28 (.A(c0nm_v0m_state_queuelen_0_), .B(c0nm_v0m_n17), .C(c0nm_v0m_state_queuelen_1_), .Y(c0nm_v0m_n14));
  // BSIM@ modules: mx16 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0nm_v0m_u16 (.A(c0nm_v0m_state_queuelen_0_), .B(c0nm_v0m_n18), .S0(c0nm_v0m_state_queuelen_1_), .Y(c0nm_v0m_n15));
  AOI21_X0P5M_A12TR c0nm_v0m_u20 (.A0(c0nm_v0m_n23), .A1(c0nm_v0m_n22), .B0(c0nm_v0m_n24), .Y(c0nm_v0m_n16));
  INV_X0P5B_A12TR c0nm_v0m_u29 (.A(c0nm_v0m_state_queuelen_2_), .Y(c0nm_v0m_n17));
  NAND3_X0P5A_A12TR c0nm_v0m_u27 (.A(c0nm_v0m_n14), .B(c0nm_v0m_n9), .C(c0nm_n2), .Y(c0nm_v0m_n18));
  // BSIM@ modules: mx16 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0nm_v0m_u18 (.A(c0nm_v0m_n20), .B(c0nm_v0m_n21), .S0(c0nm_v0m_state_queuelen_1_), .Y(c0nm_v0m_n19));
  // BSIM@ modules: mx15 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0nm_v0m_u4 (.A(c0nm_v0m_n3), .B(c0nm_routewire[1]), .S0(c0nm_v0m_n4), .Y(c0nm_v0m_n2));
  MXIT2_X0P5M_A12TR c0nm_v0m_u21 (.A(c0nm_v0m_n18), .B(c0nm_v0m_n25), .S0(c0nm_v0m_n23), .Y(c0nm_v0m_n20));
  OAI21_X0P5M_A12TR c0nm_v0m_u19 (.A0(c0nm_v0m_n22), .A1(c0nm_v0m_n23), .B0(c0nm_v0m_n16), .Y(c0nm_v0m_n21));
  INV_X0P5B_A12TR c0nm_v0m_u26 (.A(c0nm_v0m_n18), .Y(c0nm_v0m_n22));
  INV_X0P5B_A12TR c0nm_v0m_u34 (.A(c0nm_v0m_state_queuelen_0_), .Y(c0nm_v0m_n23));
  AOI21_X0P5M_A12TR c0nm_v0m_u25 (.A0(c0nm_v0m_n26), .A1(c0nm_v0m_n13), .B0(c0nm_v0m_n22), .Y(c0nm_v0m_n24));
  NAND2_X0P5A_A12TR c0nm_v0m_u22 (.A(c0nm_v0m_n13), .B(c0nm_v0m_n26), .Y(c0nm_v0m_n25));
  INV_X0P5B_A12TR c0nm_v0m_u33 (.A(c0nm_v0m_full), .Y(c0nm_v0m_n26));
  XNOR2_X0P5M_A12TR c0nm_v0m_u24 (.A(c0nm_v0m_n23), .B(c0nm_v0m_n24), .Y(c0nm_v0m_n27));
  OAI31_X0P5M_A12TR c0nm_v0m_u32 (.A0(c0nm_v0m_n29), .A1(tailout_0), .A2(c0nm_v0m_state_status_0_), .B0(c0nm_v0m_n5), .Y(c0nm_v0m_n28));
  INV_X0P5B_A12TR c0nm_v0m_u40 (.A(c0nm_v0m_state_status_1_), .Y(c0nm_v0m_n29));
  // BSIM@ modules: mx324 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_v0m_u5 (.A(swalloc_req_0[1]), .B(c0nm_v0m_n5), .Y(c0nm_v0m_n3));
  // BSIM@ modules: mx358 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0nm_v0m_u6 (.A(c0nm_v0m_n1), .B(c0nm_v0m_n6), .Y(c0nm_v0m_n30));
  // BSIM@ modules: mx358 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0nm_v0m_u3 (.A(c0nm_v0m_n1), .B(c0nm_v0m_n2), .Y(c0nm_v0m_n31));
  OA211_X0P5M_A12TR c0nm_v0m_u36 (.A0(c0nm_routewire[1]), .A1(c0nm_routewire[0]), .B0(c0nm_v0m_state_status_0_), .C0(c0nm_v0m_state_status_1_), .Y(c0nm_v0m_n4));
  OAI211_X0P5M_A12TR c0nm_v0m_u39 (.A0(swalloc_resp_0[1]), .A1(swalloc_resp_0[0]), .B0(c0nm_v0m_n29), .C0(c0nm_v0m_state_status_0_), .Y(c0nm_v0m_n5));
  AO1B2_X0P5M_A12TR c0nm_v0m_u37 (.A0N(c0nm_v0m_n8), .B0(c0nm_v0m_n5), .B1(c0nm_v0m_state_status_0_), .Y(c0nm_v0m_n57));
  AO21A1AI2_X0P5M_A12TR c0nm_v0m_u35 (.A0(c0nm_v0m_n29), .A1(c0nm_v0m_n5), .B0(c0nm_v0m_n4), .C0(c0nm_v0m_n8), .Y(c0nm_v0m_n58));
  // BSIM@ modules: mx15 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0nm_v0m_u7 (.A(c0nm_v0m_n7), .B(c0nm_routewire[0]), .S0(c0nm_v0m_n4), .Y(c0nm_v0m_n6));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0nm_v0m_u23 (.A(reset), .B(c0nm_v0m_n27), .Y(c0nm_v0m_n61));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0nm_v0m_u17 (.A(reset), .B(c0nm_v0m_n19), .Y(c0nm_v0m_n62));
  AOI211_X0P5M_A12TR c0nm_v0m_u15 (.A0(c0nm_v0m_n15), .A1(c0nm_v0m_n16), .B0(c0nm_v0m_n17), .C0(reset), .Y(c0nm_v0m_n63));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0nm_v0m_u11 (.A(reset), .B(c0nm_v0m_n10), .Y(c0nm_v0m_n64));
  // BSIM@ modules: mx325 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_v0m_u8 (.A(swalloc_req_0[0]), .B(c0nm_v0m_n5), .Y(c0nm_v0m_n7));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0nm_v0m_u38 (.A(reset), .B(tailout_0), .Y(c0nm_v0m_n8));
  OAI31_X0P5M_A12TR c0nm_v0m_u31 (.A0(c0nm_v0m_state_queuelen_0_), .A1(c0nm_v0m_state_queuelen_2_), .A2(c0nm_v0m_state_queuelen_1_), .B0(c0nm_v0m_n28), .Y(c0nm_v0m_n9));
  DFFQ_X1M_A12TR c0nm_v0m_state_queuelen_reg_0_ (.CK(clk), .Q(c0nm_v0m_state_queuelen_0_), .D(c0nm_v0m_n61));
  DFFQ_X1M_A12TR c0nm_v0m_state_queuelen_reg_1_ (.CK(clk), .Q(c0nm_v0m_state_queuelen_1_), .D(c0nm_v0m_n62));
  DFFQ_X1M_A12TR c0nm_v0m_state_queuelen_reg_2_ (.CK(clk), .Q(c0nm_v0m_state_queuelen_2_), .D(c0nm_v0m_n63));
  DFFQ_X1M_A12TR c0nm_v0m_state_status_reg_0_ (.CK(clk), .Q(c0nm_v0m_state_status_0_), .D(c0nm_v0m_n57));
  DFFQ_X1M_A12TR c0nm_v0m_state_status_reg_1_ (.CK(clk), .Q(c0nm_v0m_state_status_1_), .D(c0nm_v0m_n58));
  TIELO_X1M_A12TR c0sm_u2 (.Y(c0sm__logic0_));
  TIELO_X1M_A12TR c0sm_b0m_u3 (.Y(c0sm_b0m__logic0_));
  DFFQ_X1M_A12TR c0sm_b0m_dqenablereg_reg (.CK(clk), .Q(c0sm_b0m_dqenablereg), .D(c0sm_b0m_n9));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u255 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n180), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n71), .C0(c0sm_b0m_v0m_n274), .Y(c0sm_b0m_headflit_10_));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u250 (.A0(c0sm_b0m_v0m_n186), .A1(c0sm_b0m_v0m_n187), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n21), .C0(c0sm_b0m_v0m_n273), .Y(c0sm_b0m_headflit_11_));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u215 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n168), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n65), .C0(c0sm_b0m_v0m_n266), .Y(c0sm_b0m_headflit_8_));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u210 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n174), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n68), .C0(c0sm_b0m_v0m_n265), .Y(c0sm_b0m_headflit_9_));
  // BSIM@ modules: mx345 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR c0sm_b0m_u14 (.A(flitin_1[1]), .B(flitin_1[0]), .Y(c0sm_b0m_n2));
  // BSIM@ modules: mx361 
  // BSIM@ covered_modules=1 :   NOR2B_X0P5M_A12TR c0sm_b0m_u27 (.AN(debitout_1), .B(reset), .Y(c0sm_b0m_n9));
  // BSIM@ modules: mx246 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_0_ (.CK(clk), .Q(c0sm_b0m_rdata[0]), .D(c0sm_b0m_v0m_n331));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_10_ (.CK(clk), .Q(c0sm_b0m_rdata[10]), .D(c0sm_b0m_v0m_n341));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_11_ (.CK(clk), .Q(c0sm_b0m_rdata[11]), .D(c0sm_b0m_v0m_n342));
  // BSIM@ modules: mx246 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_1_ (.CK(clk), .Q(c0sm_b0m_rdata[1]), .D(c0sm_b0m_v0m_n332));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_2_ (.CK(clk), .Q(c0sm_b0m_rdata[2]), .D(c0sm_b0m_v0m_n333));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_3_ (.CK(clk), .Q(c0sm_b0m_rdata[3]), .D(c0sm_b0m_v0m_n334));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_4_ (.CK(clk), .Q(c0sm_b0m_rdata[4]), .D(c0sm_b0m_v0m_n335));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_5_ (.CK(clk), .Q(c0sm_b0m_rdata[5]), .D(c0sm_b0m_v0m_n336));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_6_ (.CK(clk), .Q(c0sm_b0m_rdata[6]), .D(c0sm_b0m_v0m_n337));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_7_ (.CK(clk), .Q(c0sm_b0m_rdata[7]), .D(c0sm_b0m_v0m_n338));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_8_ (.CK(clk), .Q(c0sm_b0m_rdata[8]), .D(c0sm_b0m_v0m_n339));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_9_ (.CK(clk), .Q(c0sm_b0m_rdata[9]), .D(c0sm_b0m_v0m_n340));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_0_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers0_0_), .D(c0sm_b0m_v0m_n295));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_10_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers0_10_), .D(c0sm_b0m_v0m_n305));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_11_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers0_11_), .D(c0sm_b0m_v0m_n306));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_1_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers0_1_), .D(c0sm_b0m_v0m_n296));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_2_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers0_2_), .D(c0sm_b0m_v0m_n297));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_3_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers0_3_), .D(c0sm_b0m_v0m_n298));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_4_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers0_4_), .D(c0sm_b0m_v0m_n299));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_5_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers0_5_), .D(c0sm_b0m_v0m_n300));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_6_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers0_6_), .D(c0sm_b0m_v0m_n301));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_7_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers0_7_), .D(c0sm_b0m_v0m_n302));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_8_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers0_8_), .D(c0sm_b0m_v0m_n303));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers0_reg_9_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers0_9_), .D(c0sm_b0m_v0m_n304));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_0_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers2_0_), .D(c0sm_b0m_v0m_n319));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_10_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers2_10_), .D(c0sm_b0m_v0m_n329));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_11_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers2_11_), .D(c0sm_b0m_v0m_n330));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_1_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers2_1_), .D(c0sm_b0m_v0m_n320));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_2_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers2_2_), .D(c0sm_b0m_v0m_n321));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_3_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers2_3_), .D(c0sm_b0m_v0m_n322));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_4_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers2_4_), .D(c0sm_b0m_v0m_n323));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_5_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers2_5_), .D(c0sm_b0m_v0m_n324));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_6_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers2_6_), .D(c0sm_b0m_v0m_n325));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_7_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers2_7_), .D(c0sm_b0m_v0m_n326));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_8_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers2_8_), .D(c0sm_b0m_v0m_n327));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers2_reg_9_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers2_9_), .D(c0sm_b0m_v0m_n328));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_0_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers3_0_), .D(c0sm_b0m_v0m_n284));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_10_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers3_10_), .D(c0sm_b0m_v0m_n294));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_11_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers3_11_), .D(c0sm_b0m_v0m_n283));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_1_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers3_1_), .D(c0sm_b0m_v0m_n285));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_2_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers3_2_), .D(c0sm_b0m_v0m_n286));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_3_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers3_3_), .D(c0sm_b0m_v0m_n287));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_4_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers3_4_), .D(c0sm_b0m_v0m_n288));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_5_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers3_5_), .D(c0sm_b0m_v0m_n289));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_6_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers3_6_), .D(c0sm_b0m_v0m_n290));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_7_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers3_7_), .D(c0sm_b0m_v0m_n291));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_8_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers3_8_), .D(c0sm_b0m_v0m_n292));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_buffers3_reg_9_ (.CK(clk), .Q(c0sm_b0m_v0m_buffers3_9_), .D(c0sm_b0m_v0m_n293));
  // BSIM@ modules: mx406 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0sm_b0m_v0m_head_reg_0_ (.CK(clk), .Q(c0sm_b0m_v0m_head_0_), .D(c0sm_b0m_v0m_n280));
  // BSIM@ modules: mx406 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0sm_b0m_v0m_head_reg_1_ (.CK(clk), .Q(c0sm_b0m_v0m_head_1_), .D(c0sm_b0m_v0m_n281));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_head_reg_2_ (.CK(clk), .Q(c0sm_b0m_v0m_head_2_), .D(c0sm_b0m_v0m_n282));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u7 (.A(c0sm_b0m_v0m_n8), .Y(c0sm_b0m_v0m_n1));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0sm_b0m_v0m_u208 (.A(c0sm_b0m_v0m_n11), .B(reset), .Y(c0sm_b0m_v0m_n10));
  // BSIM@ modules: mx281 
  // BSIM@ covered_modules=1 :   NAND3_X0P5A_A12TR c0sm_b0m_v0m_u80 (.A(c0sm_b0m_v0m_n95), .B(c0sm_b0m_v0m_n94), .C(c0sm_b0m_v0m_n72), .Y(c0sm_b0m_v0m_n100));
  // BSIM@ modules: mx132 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0sm_b0m_v0m_u68 (.A0(c0sm_b0m_v0m_n99), .A1(c0sm_b0m_v0m_n31), .B0(c0sm_b0m_v0m_n100), .B1(c0sm_b0m_v0m_n32), .C0(reset), .Y(c0sm_b0m_v0m_n101));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR c0sm_b0m_v0m_u82 (.A(c0sm_b0m_v0m_n99), .B(c0nm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n102));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u79 (.A(c0sm_b0m_v0m_n98), .B(c0nm_b0m_v0m_n4), .C(c0sm_b0m_v0m_n100), .Y(c0sm_b0m_v0m_n103));
  // BSIM@ modules: mx316 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u176 (.A(c0sm_b0m_v0m_n192), .Y(c0sm_b0m_v0m_n104));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u275 (.A(c0sm_b0m_v0m_buffers2_0_), .Y(c0sm_b0m_v0m_n105));
  // BSIM@ modules: mx370 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0sm_b0m_v0m_u85 (.A0(c0sm_b0m_v0m_n108), .A1(c0sm_b0m_v0m_n25), .B0(c0sm_b0m_v0m_n109), .B1(c0sm_b0m_v0m_n27), .C0(reset), .Y(c0sm_b0m_v0m_n106));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u167 (.A(c0sm_b0m_v0m_n187), .B(c0nm_b0m_v0m_n4), .C(c0sm_b0m_v0m_n94), .Y(c0sm_b0m_v0m_n107));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u179 (.A(c0sm_b0m_v0m_n94), .Y(c0sm_b0m_v0m_n108));
  // BSIM@ modules: mx281 
  // BSIM@ covered_modules=1 :   NAND3_X0P5A_A12TR c0sm_b0m_v0m_u164 (.A(c0sm_b0m_v0m_n93), .B(c0sm_b0m_v0m_n95), .C(c0sm_b0m_v0m_n72), .Y(c0sm_b0m_v0m_n109));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0sm_b0m_v0m_u209 (.A(debitout_1), .B(reset), .Y(c0sm_b0m_v0m_n11));
  // BSIM@ modules: mx316 
  // BSIM@ covered_modules=1 :   OR2_X0P5M_A12TR c0sm_b0m_v0m_u173 (.A(c0sm_b0m_v0m_n187), .B(debitout_1), .Y(c0sm_b0m_v0m_n110));
  NAND4_X0P5A_A12TR c0sm_b0m_v0m_u174 (.A(c0sm_b0m_v0m_n96), .B(c0sm_b0m_v0m_n104), .C(c0sm_b0m_v0m_n187), .D(c0sm_v0m_n9), .Y(c0sm_b0m_v0m_n111));
  // BSIM@ modules: mx194 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0sm_b0m_v0m_u87 (.A0(c0sm_b0m_v0m_n113), .A1(c0sm_b0m_v0m_n114), .B0(c0sm_b0m_v0m_buffers0_0_), .B1(c0sm_b0m_v0m_n115), .C0(debitout_1), .Y(c0sm_b0m_v0m_n112));
  // BSIM@ modules: mx316 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0sm_b0m_v0m_u171 (.A(c0sm_b0m_v0m_n104), .B(debitout_1), .Y(c0sm_b0m_v0m_n113));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u270 (.A(c0sm_b0m_v0m_n343), .Y(c0sm_b0m_v0m_n114));
  // BSIM@ modules: mx316 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0sm_b0m_v0m_u172 (.A(c0sm_b0m_v0m_n96), .B(debitout_1), .Y(c0sm_b0m_v0m_n115));
  // BSIM@ modules: mx338 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u98 (.A(c0sm_b0m_v0m_n128), .Y(c0sm_b0m_v0m_n116));
  // BSIM@ modules: mx88 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u90 (.A0(c0sm_b0m_v0m_buffers0_0_), .A1(c0sm_b0m_v0m_n120), .B0(c0sm_b0m_v0m_buffers2_0_), .B1(c0sm_b0m_v0m_n121), .Y(c0sm_b0m_v0m_n117));
  // BSIM@ modules: mx65 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u89 (.A0(c0sm_b0m_v0m_n119), .A1(c0sm_b0m_v0m_n114), .B0(flitin_1[0]), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n118));
  // BSIM@ modules: mx338 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0sm_b0m_v0m_u191 (.A(c0sm_b0m_v0m_n93), .B(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n119));
  AOI21_X0P5M_A12TR c0sm_b0m_v0m_u16 (.A0(c0nm_b0m_v0m_n4), .A1(c0sm_b0m_v0m_n16), .B0(c0sm_b0m_v0m_n11), .Y(c0sm_b0m_v0m_n12));
  // BSIM@ modules: mx359 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0sm_b0m_v0m_u185 (.A(c0sm_b0m_v0m_n95), .B(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n120));
  // BSIM@ modules: mx359 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0sm_b0m_v0m_u187 (.A(c0sm_b0m_v0m_n94), .B(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n121));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u267 (.A(c0sm_b0m_v0m_buffers2_1_), .Y(c0sm_b0m_v0m_n122));
  // BSIM@ modules: mx370 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0sm_b0m_v0m_u92 (.A0(c0sm_b0m_v0m_n108), .A1(c0sm_b0m_v0m_n31), .B0(c0sm_b0m_v0m_n109), .B1(c0sm_b0m_v0m_n32), .C0(reset), .Y(c0sm_b0m_v0m_n123));
  // BSIM@ modules: mx194 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0sm_b0m_v0m_u94 (.A0(c0sm_b0m_v0m_n113), .A1(c0sm_b0m_v0m_n125), .B0(c0sm_b0m_v0m_buffers0_1_), .B1(c0sm_b0m_v0m_n115), .C0(debitout_1), .Y(c0sm_b0m_v0m_n124));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u265 (.A(c0sm_b0m_v0m_n344), .Y(c0sm_b0m_v0m_n125));
  // BSIM@ modules: mx88 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u97 (.A0(c0sm_b0m_v0m_buffers0_1_), .A1(c0sm_b0m_v0m_n120), .B0(c0sm_b0m_v0m_buffers2_1_), .B1(c0sm_b0m_v0m_n121), .Y(c0sm_b0m_v0m_n126));
  // BSIM@ modules: mx65 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u96 (.A0(c0sm_b0m_v0m_n119), .A1(c0sm_b0m_v0m_n125), .B0(flitin_1[1]), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n127));
  // BSIM@ modules: mx338 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0sm_b0m_v0m_u182 (.A(c0sm_b0m_v0m_n28), .B(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n128));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR c0sm_b0m_v0m_u178 (.A(c0sm_b0m_v0m_n108), .B(c0nm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n129));
  NAND2_X0P5A_A12TR c0sm_b0m_v0m_u14 (.A(c0sm_b0m_v0m_n10), .B(c0sm_b0m_v0m_head_0_), .Y(c0sm_b0m_v0m_n13));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u163 (.A(c0sm_b0m_v0m_n107), .B(c0nm_b0m_v0m_n4), .C(c0sm_b0m_v0m_n109), .Y(c0sm_b0m_v0m_n130));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u249 (.A(c0sm_b0m_v0m_buffers2_2_), .Y(c0sm_b0m_v0m_n131));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u101 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n35), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n131), .C0(c0sm_b0m_v0m_n133), .Y(c0sm_b0m_v0m_n132));
  // BSIM@ modules: mx99 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u102 (.A0(c0sm_b0m_v0m_buffers0_2_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n134), .Y(c0sm_b0m_v0m_n133));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u247 (.A(c0sm_b0m_v0m_n345), .Y(c0sm_b0m_v0m_n134));
  // BSIM@ modules: mx338 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u190 (.A(c0sm_b0m_v0m_n119), .Y(c0sm_b0m_v0m_n135));
  // BSIM@ modules: mx88 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u105 (.A0(c0sm_b0m_v0m_buffers2_2_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_2_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n136));
  // BSIM@ modules: mx66 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u104 (.A0(c0sm_b0m_v0m_buffers3_2_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_2_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n137));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u244 (.A(c0sm_b0m_v0m_buffers2_3_), .Y(c0sm_b0m_v0m_n138));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u108 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n38), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n138), .C0(c0sm_b0m_v0m_n140), .Y(c0sm_b0m_v0m_n139));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u13 (.A(c0sm_b0m_v0m_head_1_), .Y(c0sm_b0m_v0m_n14));
  // BSIM@ modules: mx99 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u109 (.A0(c0sm_b0m_v0m_buffers0_3_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n141), .Y(c0sm_b0m_v0m_n140));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u242 (.A(c0sm_b0m_v0m_n346), .Y(c0sm_b0m_v0m_n141));
  // BSIM@ modules: mx88 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u112 (.A0(c0sm_b0m_v0m_buffers2_3_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_3_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n142));
  // BSIM@ modules: mx66 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u111 (.A0(c0sm_b0m_v0m_buffers3_3_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_3_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n143));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u239 (.A(c0sm_b0m_v0m_buffers2_4_), .Y(c0sm_b0m_v0m_n144));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u115 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n41), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n144), .C0(c0sm_b0m_v0m_n146), .Y(c0sm_b0m_v0m_n145));
  // BSIM@ modules: mx99 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u116 (.A0(c0sm_b0m_v0m_buffers0_4_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n147), .Y(c0sm_b0m_v0m_n146));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u237 (.A(c0sm_b0m_v0m_n347), .Y(c0sm_b0m_v0m_n147));
  // BSIM@ modules: mx88 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u119 (.A0(c0sm_b0m_v0m_buffers2_4_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_4_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n148));
  // BSIM@ modules: mx66 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u118 (.A0(c0sm_b0m_v0m_buffers3_4_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_4_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n149));
  // BSIM@ modules: mx316 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u277 (.A(c0sm_b0m_v0m_head_2_), .Y(c0sm_b0m_v0m_n15));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u234 (.A(c0sm_b0m_v0m_buffers2_5_), .Y(c0sm_b0m_v0m_n150));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u122 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n44), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n150), .C0(c0sm_b0m_v0m_n152), .Y(c0sm_b0m_v0m_n151));
  // BSIM@ modules: mx99 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u123 (.A0(c0sm_b0m_v0m_buffers0_5_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n153), .Y(c0sm_b0m_v0m_n152));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u232 (.A(c0sm_b0m_v0m_n348), .Y(c0sm_b0m_v0m_n153));
  // BSIM@ modules: mx88 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u126 (.A0(c0sm_b0m_v0m_buffers2_5_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_5_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n154));
  // BSIM@ modules: mx66 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u125 (.A0(c0sm_b0m_v0m_buffers3_5_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_5_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n155));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u229 (.A(c0sm_b0m_v0m_buffers2_6_), .Y(c0sm_b0m_v0m_n156));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u129 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n47), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n156), .C0(c0sm_b0m_v0m_n158), .Y(c0sm_b0m_v0m_n157));
  // BSIM@ modules: mx99 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u130 (.A0(c0sm_b0m_v0m_buffers0_6_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n159), .Y(c0sm_b0m_v0m_n158));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u227 (.A(c0sm_b0m_v0m_n349), .Y(c0sm_b0m_v0m_n159));
  // BSIM@ modules: mx316 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u278 (.A(c0sm_b0m_v0m_head_0_), .Y(c0sm_b0m_v0m_n16));
  // BSIM@ modules: mx88 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u133 (.A0(c0sm_b0m_v0m_buffers2_6_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_6_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n160));
  // BSIM@ modules: mx66 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u132 (.A0(c0sm_b0m_v0m_buffers3_6_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_6_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n161));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u224 (.A(c0sm_b0m_v0m_buffers2_7_), .Y(c0sm_b0m_v0m_n162));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u136 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n62), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n162), .C0(c0sm_b0m_v0m_n164), .Y(c0sm_b0m_v0m_n163));
  // BSIM@ modules: mx99 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u137 (.A0(c0sm_b0m_v0m_buffers0_7_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n165), .Y(c0sm_b0m_v0m_n164));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u222 (.A(c0sm_b0m_v0m_n350), .Y(c0sm_b0m_v0m_n165));
  // BSIM@ modules: mx88 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u140 (.A0(c0sm_b0m_v0m_buffers2_7_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_7_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n166));
  // BSIM@ modules: mx66 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u139 (.A0(c0sm_b0m_v0m_buffers3_7_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_7_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n167));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u219 (.A(c0sm_b0m_v0m_buffers2_8_), .Y(c0sm_b0m_v0m_n168));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u143 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n65), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n168), .C0(c0sm_b0m_v0m_n170), .Y(c0sm_b0m_v0m_n169));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u168 (.A(c0sm_b0m_v0m_n188), .Y(c0sm_b0m_v0m_n17));
  // BSIM@ modules: mx99 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u144 (.A0(c0sm_b0m_v0m_buffers0_8_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n171), .Y(c0sm_b0m_v0m_n170));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u217 (.A(c0sm_b0m_v0m_n351), .Y(c0sm_b0m_v0m_n171));
  AND4_X0P5M_A12TR c0sm_b0m_v0m_u260 (.A(debitout_1), .B(c0sm_headflit[0]), .C(c0sm_b0m_v0m_n264), .D(c0nm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n1710));
  // BSIM@ modules: mx88 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u147 (.A0(c0sm_b0m_v0m_buffers2_8_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_8_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n172));
  // BSIM@ modules: mx66 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u146 (.A0(c0sm_b0m_v0m_buffers3_8_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_8_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n173));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u214 (.A(c0sm_b0m_v0m_buffers2_9_), .Y(c0sm_b0m_v0m_n174));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u150 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n68), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n174), .C0(c0sm_b0m_v0m_n176), .Y(c0sm_b0m_v0m_n175));
  // BSIM@ modules: mx99 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u151 (.A0(c0sm_b0m_v0m_buffers0_9_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n177), .Y(c0sm_b0m_v0m_n176));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u212 (.A(c0sm_b0m_v0m_n352), .Y(c0sm_b0m_v0m_n177));
  // BSIM@ modules: mx88 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u154 (.A0(c0sm_b0m_v0m_buffers2_9_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_9_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n178));
  // BSIM@ modules: mx66 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u153 (.A0(c0sm_b0m_v0m_buffers3_9_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_9_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n179));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u32 (.A(c0sm_b0m_v0m_n22), .B(c0nm_b0m_v0m_n4), .C(c0sm_b0m_v0m_n28), .Y(c0sm_b0m_v0m_n18));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u259 (.A(c0sm_b0m_v0m_buffers2_10_), .Y(c0sm_b0m_v0m_n180));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u157 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n71), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n180), .C0(c0sm_b0m_v0m_n182), .Y(c0sm_b0m_v0m_n181));
  // BSIM@ modules: mx99 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u158 (.A0(c0sm_b0m_v0m_buffers0_10_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n183), .Y(c0sm_b0m_v0m_n182));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u257 (.A(c0sm_b0m_v0m_n353), .Y(c0sm_b0m_v0m_n183));
  // BSIM@ modules: mx88 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u161 (.A0(c0sm_b0m_v0m_buffers2_10_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_10_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n184));
  // BSIM@ modules: mx66 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u160 (.A0(c0sm_b0m_v0m_buffers3_10_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_10_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n185));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u254 (.A(c0sm_b0m_v0m_buffers2_11_), .Y(c0sm_b0m_v0m_n186));
  // BSIM@ modules: mx316 
  // BSIM@ covered_modules=1 :   NAND3_X0P5A_A12TR c0sm_b0m_v0m_u276 (.A(c0sm_b0m_v0m_n16), .B(c0sm_b0m_v0m_n15), .C(c0sm_b0m_v0m_head_1_), .Y(c0sm_b0m_v0m_n187));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u169 (.A0(c0sm_b0m_v0m_n21), .A1(c0sm_b0m_v0m_n111), .B0(c0sm_b0m_v0m_n186), .B1(c0sm_b0m_v0m_n110), .C0(c0sm_b0m_v0m_n189), .Y(c0sm_b0m_v0m_n188));
  // BSIM@ modules: mx99 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u170 (.A0(c0sm_b0m_v0m_n115), .A1(c0sm_b0m_v0m_buffers0_11_), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n190), .Y(c0sm_b0m_v0m_n189));
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u180 (.A0(c0sm_b0m_v0m_n354), .A1(c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n194), .C0(c0sm_b0m_v0m_n195), .Y(c0sm_b0m_v0m_n19));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u252 (.A(c0sm_b0m_v0m_n354), .Y(c0sm_b0m_v0m_n190));
  // BSIM@ modules: mx316 
  // BSIM@ covered_modules=1 :   NOR3_X0P5A_A12TR c0sm_b0m_v0m_u271 (.A(c0sm_b0m_v0m_head_1_), .B(c0sm_b0m_v0m_head_2_), .C(c0sm_b0m_v0m_n16), .Y(c0sm_b0m_v0m_n192));
  // BSIM@ modules: mx316 
  // BSIM@ covered_modules=1 :   NOR3_X0P5A_A12TR c0sm_b0m_v0m_u272 (.A(c0sm_b0m_v0m_head_1_), .B(c0sm_b0m_v0m_head_2_), .C(c0sm_b0m_v0m_head_0_), .Y(c0sm_b0m_v0m_n193));
  // BSIM@ modules: mx88 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u184 (.A0(c0sm_b0m_v0m_buffers2_11_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_11_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n194));
  // BSIM@ modules: mx66 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u181 (.A0(c0sm_b0m_v0m_buffers3_11_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_n2), .B1(c0sm_b0m_wdata_11_), .Y(c0sm_b0m_v0m_n195));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR c0sm_b0m_v0m_u4 (.A(c0sm_b0m_v0m_n1), .B(c0nm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n2));
  // BSIM@ modules: mx346 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR c0sm_b0m_v0m_u31 (.A(c0sm_b0m_v0m_n26), .B(c0nm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n20));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u253 (.A(c0sm_b0m_v0m_buffers3_11_), .Y(c0sm_b0m_v0m_n21));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u33 (.A(c0sm_b0m_v0m_n72), .B(c0nm_b0m_v0m_n4), .C(c0sm_b0m_v0m_n73), .Y(c0sm_b0m_v0m_n22));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u273 (.A(c0sm_b0m_v0m_buffers3_0_), .Y(c0sm_b0m_v0m_n23));
  // BSIM@ modules: mx373 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0sm_b0m_v0m_u19 (.A0(c0sm_b0m_v0m_n25), .A1(c0sm_b0m_v0m_n26), .B0(c0sm_b0m_v0m_n27), .B1(c0sm_b0m_v0m_n28), .C0(reset), .Y(c0sm_b0m_v0m_n24));
  OAI211_X0P5M_A12TR c0sm_b0m_v0m_u88 (.A0(c0sm_b0m_v0m_n116), .A1(c0sm_b0m_v0m_n23), .B0(c0sm_b0m_v0m_n117), .C0(c0sm_b0m_v0m_n118), .Y(c0sm_b0m_v0m_n25));
  // BSIM@ modules: mx281 
  // BSIM@ covered_modules=1 :   OAI21_X0P5M_A12TR c0sm_b0m_v0m_u166 (.A0(c0sm_b0m_v0m_n3), .A1(c0sm_b0m_v0m_n7), .B0(c0sm_b0m_v0m_n355), .Y(c0sm_b0m_v0m_n26));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   NAND2B_X0P5M_A12TR c0sm_b0m_v0m_u195 (.AN(c0sm_headflit[0]), .B(c0nm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n262));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR c0sm_b0m_v0m_u197 (.A(c0sm_b0m_v0m_n264), .B(c0nm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n263));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u262 (.A(c0sm_headflit[1]), .Y(c0sm_b0m_v0m_n264));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u211 (.A0(c0sm_b0m_v0m_buffers0_9_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n177), .Y(c0sm_b0m_v0m_n265));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u216 (.A0(c0sm_b0m_v0m_buffers0_8_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n171), .Y(c0sm_b0m_v0m_n266));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u221 (.A0(c0sm_b0m_v0m_buffers0_7_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n165), .Y(c0sm_b0m_v0m_n267));
  // BSIM@ modules: mx77 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u226 (.A0(c0sm_b0m_v0m_buffers0_6_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n159), .Y(c0sm_b0m_v0m_n268));
  // BSIM@ modules: mx77 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u231 (.A0(c0sm_b0m_v0m_buffers0_5_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n153), .Y(c0sm_b0m_v0m_n269));
  // BSIM@ modules: mx244 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u86 (.A0(c0sm_b0m_v0m_n110), .A1(c0sm_b0m_v0m_n105), .B0(c0sm_b0m_v0m_n111), .B1(c0sm_b0m_v0m_n23), .C0(c0sm_b0m_v0m_n112), .Y(c0sm_b0m_v0m_n27));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u236 (.A0(c0sm_b0m_v0m_buffers0_4_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n147), .Y(c0sm_b0m_v0m_n270));
  // BSIM@ modules: mx77 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u241 (.A0(c0sm_b0m_v0m_buffers0_3_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n141), .Y(c0sm_b0m_v0m_n271));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u246 (.A0(c0sm_b0m_v0m_buffers0_2_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n134), .Y(c0sm_b0m_v0m_n272));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u251 (.A0(c0sm_b0m_v0m_n193), .A1(c0sm_b0m_v0m_buffers0_11_), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n190), .Y(c0sm_b0m_v0m_n273));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u256 (.A0(c0sm_b0m_v0m_buffers0_10_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n183), .Y(c0sm_b0m_v0m_n274));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u264 (.A0(c0sm_b0m_v0m_buffers0_1_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n125), .Y(c0sm_b0m_v0m_n275));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_b0m_v0m_u269 (.A0(c0sm_b0m_v0m_buffers0_0_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n114), .Y(c0sm_b0m_v0m_n276));
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u3 (.A(c0sm_b0m_v0m_n1), .B(c0sm_b0m_v0m_n2), .S0(c0sm_b0m_v0m_n3), .Y(c0sm_b0m_v0m_n277));
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u5 (.A(c0sm_b0m_v0m_n5), .B(c0sm_b0m_v0m_n6), .S0(c0sm_b0m_v0m_n7), .Y(c0sm_b0m_v0m_n278));
  OA21A1OI2_X0P5M_A12TR c0sm_b0m_v0m_u8 (.A0(c0sm_b0m_v0m_tail_1_), .A1(reset), .B0(c0sm_b0m_v0m_n5), .C0(c0sm_b0m_v0m_n355), .Y(c0sm_b0m_v0m_n279));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u183 (.A(c0sm_b0m_v0m_n95), .B(c0sm_b0m_v0m_n94), .C(c0sm_b0m_v0m_n93), .Y(c0sm_b0m_v0m_n28));
  MXT2_X0P5M_A12TR c0sm_b0m_v0m_u11 (.A(c0sm_b0m_v0m_n10), .B(c0sm_b0m_v0m_n11), .S0(c0sm_b0m_v0m_head_0_), .Y(c0sm_b0m_v0m_n280));
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u12 (.A(c0sm_b0m_v0m_n12), .B(c0sm_b0m_v0m_n13), .S0(c0sm_b0m_v0m_n14), .Y(c0sm_b0m_v0m_n281));
  OA21A1OI2_X0P5M_A12TR c0sm_b0m_v0m_u15 (.A0(reset), .A1(c0sm_b0m_v0m_head_1_), .B0(c0sm_b0m_v0m_n12), .C0(c0sm_b0m_v0m_n15), .Y(c0sm_b0m_v0m_n282));
  // BSIM@ modules: mx109 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u17 (.A0(c0sm_b0m_v0m_n17), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n19), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n21), .C1(c0sm_b0m_v0m_n22), .Y(c0sm_b0m_v0m_n283));
  // BSIM@ modules: mx373 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u18 (.A(c0sm_b0m_v0m_n23), .B(c0sm_b0m_v0m_n24), .S0(c0sm_b0m_v0m_n22), .Y(c0sm_b0m_v0m_n284));
  // BSIM@ modules: mx373 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u20 (.A(c0sm_b0m_v0m_n29), .B(c0sm_b0m_v0m_n30), .S0(c0sm_b0m_v0m_n22), .Y(c0sm_b0m_v0m_n285));
  // BSIM@ modules: mx109 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u22 (.A0(c0sm_b0m_v0m_n33), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n34), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n35), .Y(c0sm_b0m_v0m_n286));
  // BSIM@ modules: mx109 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u23 (.A0(c0sm_b0m_v0m_n36), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n37), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n38), .Y(c0sm_b0m_v0m_n287));
  // BSIM@ modules: mx109 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u24 (.A0(c0sm_b0m_v0m_n39), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n40), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n41), .Y(c0sm_b0m_v0m_n288));
  // BSIM@ modules: mx109 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u25 (.A0(c0sm_b0m_v0m_n42), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n43), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n44), .Y(c0sm_b0m_v0m_n289));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u266 (.A(c0sm_b0m_v0m_buffers3_1_), .Y(c0sm_b0m_v0m_n29));
  // BSIM@ modules: mx109 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u26 (.A0(c0sm_b0m_v0m_n45), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n46), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n47), .Y(c0sm_b0m_v0m_n290));
  // BSIM@ modules: mx109 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u27 (.A0(c0sm_b0m_v0m_n48), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n49), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n62), .Y(c0sm_b0m_v0m_n291));
  // BSIM@ modules: mx109 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u28 (.A0(c0sm_b0m_v0m_n63), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n64), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n65), .Y(c0sm_b0m_v0m_n292));
  // BSIM@ modules: mx109 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u29 (.A0(c0sm_b0m_v0m_n66), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n67), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n68), .Y(c0sm_b0m_v0m_n293));
  // BSIM@ modules: mx109 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u30 (.A0(c0sm_b0m_v0m_n69), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n70), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n71), .Y(c0sm_b0m_v0m_n294));
  // BSIM@ modules: mx372 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u34 (.A(c0sm_b0m_v0m_n74), .B(c0sm_b0m_v0m_n75), .S0(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n295));
  // BSIM@ modules: mx372 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u37 (.A(c0sm_b0m_v0m_n79), .B(c0sm_b0m_v0m_n80), .S0(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n296));
  // BSIM@ modules: mx108 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u40 (.A0(c0sm_b0m_v0m_n34), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n33), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n83), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n297));
  // BSIM@ modules: mx108 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u42 (.A0(c0sm_b0m_v0m_n37), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n36), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n84), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n298));
  // BSIM@ modules: mx108 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u44 (.A0(c0sm_b0m_v0m_n40), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n39), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n85), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n299));
  // BSIM@ modules: mx281 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u189 (.A(c0sm_b0m_v0m_tail_0_), .Y(c0sm_b0m_v0m_n3));
  // BSIM@ modules: mx373 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0sm_b0m_v0m_u21 (.A0(c0sm_b0m_v0m_n31), .A1(c0sm_b0m_v0m_n26), .B0(c0sm_b0m_v0m_n32), .B1(c0sm_b0m_v0m_n28), .C0(reset), .Y(c0sm_b0m_v0m_n30));
  // BSIM@ modules: mx108 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u46 (.A0(c0sm_b0m_v0m_n43), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n42), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n86), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n300));
  // BSIM@ modules: mx108 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u48 (.A0(c0sm_b0m_v0m_n46), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n45), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n87), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n301));
  // BSIM@ modules: mx108 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u50 (.A0(c0sm_b0m_v0m_n49), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n48), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n88), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n302));
  // BSIM@ modules: mx108 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u52 (.A0(c0sm_b0m_v0m_n64), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n63), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n89), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n303));
  // BSIM@ modules: mx108 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u54 (.A0(c0sm_b0m_v0m_n67), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n66), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n90), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n304));
  // BSIM@ modules: mx108 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u56 (.A0(c0sm_b0m_v0m_n70), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n69), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n91), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n305));
  // BSIM@ modules: mx108 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u58 (.A0(c0sm_b0m_v0m_n19), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n17), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n92), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n306));
  // BSIM@ modules: mx248 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u65 (.A(c0sm_b0m_v0m_n343), .B(c0sm_b0m_v0m_n97), .S0(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n307));
  // BSIM@ modules: mx248 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u67 (.A(c0sm_b0m_v0m_n344), .B(c0sm_b0m_v0m_n101), .S0(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n308));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u69 (.A0(c0sm_b0m_v0m_n34), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n33), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n345), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n309));
  OAI211_X0P5M_A12TR c0sm_b0m_v0m_u95 (.A0(c0sm_b0m_v0m_n116), .A1(c0sm_b0m_v0m_n29), .B0(c0sm_b0m_v0m_n126), .C0(c0sm_b0m_v0m_n127), .Y(c0sm_b0m_v0m_n31));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u70 (.A0(c0sm_b0m_v0m_n37), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n36), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n346), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n310));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u71 (.A0(c0sm_b0m_v0m_n40), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n39), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n347), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n311));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u72 (.A0(c0sm_b0m_v0m_n43), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n42), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n348), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n312));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u73 (.A0(c0sm_b0m_v0m_n46), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n45), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n349), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n313));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u74 (.A0(c0sm_b0m_v0m_n49), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n48), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n350), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n314));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u75 (.A0(c0sm_b0m_v0m_n64), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n63), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n351), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n315));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u76 (.A0(c0sm_b0m_v0m_n67), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n66), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n352), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n316));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u77 (.A0(c0sm_b0m_v0m_n70), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n69), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n353), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n317));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u78 (.A0(c0sm_b0m_v0m_n19), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n17), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n354), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n318));
  // BSIM@ modules: mx370 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u84 (.A(c0sm_b0m_v0m_n105), .B(c0sm_b0m_v0m_n106), .S0(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n319));
  // BSIM@ modules: mx244 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u93 (.A0(c0sm_b0m_v0m_n110), .A1(c0sm_b0m_v0m_n122), .B0(c0sm_b0m_v0m_n111), .B1(c0sm_b0m_v0m_n29), .C0(c0sm_b0m_v0m_n124), .Y(c0sm_b0m_v0m_n32));
  // BSIM@ modules: mx370 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u91 (.A(c0sm_b0m_v0m_n122), .B(c0sm_b0m_v0m_n123), .S0(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n320));
  // BSIM@ modules: mx106 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u99 (.A0(c0sm_b0m_v0m_n34), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n33), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n131), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n321));
  // BSIM@ modules: mx106 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u106 (.A0(c0sm_b0m_v0m_n37), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n36), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n138), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n322));
  // BSIM@ modules: mx106 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u113 (.A0(c0sm_b0m_v0m_n40), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n39), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n144), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n323));
  // BSIM@ modules: mx106 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u120 (.A0(c0sm_b0m_v0m_n43), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n42), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n150), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n324));
  // BSIM@ modules: mx106 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u127 (.A0(c0sm_b0m_v0m_n46), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n45), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n156), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n325));
  // BSIM@ modules: mx106 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u134 (.A0(c0sm_b0m_v0m_n49), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n48), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n162), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n326));
  // BSIM@ modules: mx106 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u141 (.A0(c0sm_b0m_v0m_n64), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n63), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n168), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n327));
  // BSIM@ modules: mx106 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u148 (.A0(c0sm_b0m_v0m_n67), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n66), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n174), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n328));
  // BSIM@ modules: mx106 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u155 (.A0(c0sm_b0m_v0m_n70), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n69), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n180), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n329));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u100 (.A(c0sm_b0m_v0m_n132), .Y(c0sm_b0m_v0m_n33));
  // BSIM@ modules: mx106 
  // BSIM@ covered_modules=1 :   OAI222_X0P5M_A12TR c0sm_b0m_v0m_u162 (.A0(c0sm_b0m_v0m_n19), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n17), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n186), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n330));
  // BSIM@ modules: mx246 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR c0sm_b0m_v0m_u194 (.A(c0sm_b0m_v0m_n262), .B(c0sm_b0m_rdata[0]), .S0(c0sm_b0m_v0m_n11), .Y(c0sm_b0m_v0m_n331));
  // BSIM@ modules: mx246 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR c0sm_b0m_v0m_u196 (.A(c0sm_b0m_v0m_n263), .B(c0sm_b0m_rdata[1]), .S0(c0sm_b0m_v0m_n11), .Y(c0sm_b0m_v0m_n332));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0sm_b0m_v0m_u198 (.A0(c0sm_b0m_rdata[2]), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit[2]), .Y(c0sm_b0m_v0m_n333));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0sm_b0m_v0m_u199 (.A0(c0sm_b0m_rdata[3]), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit[3]), .Y(c0sm_b0m_v0m_n334));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0sm_b0m_v0m_u200 (.A0(c0sm_b0m_rdata[4]), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit[4]), .Y(c0sm_b0m_v0m_n335));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0sm_b0m_v0m_u201 (.A0(c0sm_b0m_rdata[5]), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit[5]), .Y(c0sm_b0m_v0m_n336));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0sm_b0m_v0m_u202 (.A0(c0sm_b0m_rdata[6]), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit[6]), .Y(c0sm_b0m_v0m_n337));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0sm_b0m_v0m_u203 (.A0(c0sm_b0m_rdata[7]), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit[7]), .Y(c0sm_b0m_v0m_n338));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0sm_b0m_v0m_u204 (.A0(c0sm_b0m_rdata[8]), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_b0m_headflit_8_), .Y(c0sm_b0m_v0m_n339));
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u103 (.A0(c0sm_b0m_v0m_n345), .A1(c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n136), .C0(c0sm_b0m_v0m_n137), .Y(c0sm_b0m_v0m_n34));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0sm_b0m_v0m_u205 (.A0(c0sm_b0m_rdata[9]), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_b0m_headflit_9_), .Y(c0sm_b0m_v0m_n340));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0sm_b0m_v0m_u206 (.A0(c0sm_b0m_rdata[10]), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_b0m_headflit_10_), .Y(c0sm_b0m_v0m_n341));
  // BSIM@ modules: mx250 
  // BSIM@ covered_modules=1 :   AO22_X0P5M_A12TR c0sm_b0m_v0m_u207 (.A0(c0sm_b0m_rdata[11]), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_b0m_headflit_11_), .Y(c0sm_b0m_v0m_n342));
  // BSIM@ modules: mx248 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_0_ (.CK(clk), .QN(c0sm_b0m_v0m_n343), .D(c0sm_b0m_v0m_n307));
  // BSIM@ modules: mx248 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_1_ (.CK(clk), .QN(c0sm_b0m_v0m_n344), .D(c0sm_b0m_v0m_n308));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_2_ (.CK(clk), .QN(c0sm_b0m_v0m_n345), .D(c0sm_b0m_v0m_n309));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_3_ (.CK(clk), .QN(c0sm_b0m_v0m_n346), .D(c0sm_b0m_v0m_n310));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_4_ (.CK(clk), .QN(c0sm_b0m_v0m_n347), .D(c0sm_b0m_v0m_n311));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_5_ (.CK(clk), .QN(c0sm_b0m_v0m_n348), .D(c0sm_b0m_v0m_n312));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_6_ (.CK(clk), .QN(c0sm_b0m_v0m_n349), .D(c0sm_b0m_v0m_n313));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u248 (.A(c0sm_b0m_v0m_buffers3_2_), .Y(c0sm_b0m_v0m_n35));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_7_ (.CK(clk), .QN(c0sm_b0m_v0m_n350), .D(c0sm_b0m_v0m_n314));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_8_ (.CK(clk), .QN(c0sm_b0m_v0m_n351), .D(c0sm_b0m_v0m_n315));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_9_ (.CK(clk), .QN(c0sm_b0m_v0m_n352), .D(c0sm_b0m_v0m_n316));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_10_ (.CK(clk), .QN(c0sm_b0m_v0m_n353), .D(c0sm_b0m_v0m_n317));
  // BSIM@ modules: mx252 
  // BSIM@ covered_modules=1 :   DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_11_ (.CK(clk), .QN(c0sm_b0m_v0m_n354), .D(c0sm_b0m_v0m_n318));
  DFFQN_X1M_A12TR c0sm_b0m_v0m_tail_reg_2_ (.CK(clk), .QN(c0sm_b0m_v0m_n355), .D(c0sm_b0m_v0m_n279));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u107 (.A(c0sm_b0m_v0m_n139), .Y(c0sm_b0m_v0m_n36));
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u110 (.A0(c0sm_b0m_v0m_n346), .A1(c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n142), .C0(c0sm_b0m_v0m_n143), .Y(c0sm_b0m_v0m_n37));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u243 (.A(c0sm_b0m_v0m_buffers3_3_), .Y(c0sm_b0m_v0m_n38));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u114 (.A(c0sm_b0m_v0m_n145), .Y(c0sm_b0m_v0m_n39));
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u117 (.A0(c0sm_b0m_v0m_n347), .A1(c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n148), .C0(c0sm_b0m_v0m_n149), .Y(c0sm_b0m_v0m_n40));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u238 (.A(c0sm_b0m_v0m_buffers3_4_), .Y(c0sm_b0m_v0m_n41));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u121 (.A(c0sm_b0m_v0m_n151), .Y(c0sm_b0m_v0m_n42));
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u124 (.A0(c0sm_b0m_v0m_n348), .A1(c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n154), .C0(c0sm_b0m_v0m_n155), .Y(c0sm_b0m_v0m_n43));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u233 (.A(c0sm_b0m_v0m_buffers3_5_), .Y(c0sm_b0m_v0m_n44));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u128 (.A(c0sm_b0m_v0m_n157), .Y(c0sm_b0m_v0m_n45));
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u131 (.A0(c0sm_b0m_v0m_n349), .A1(c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n160), .C0(c0sm_b0m_v0m_n161), .Y(c0sm_b0m_v0m_n46));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u228 (.A(c0sm_b0m_v0m_buffers3_6_), .Y(c0sm_b0m_v0m_n47));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u135 (.A(c0sm_b0m_v0m_n163), .Y(c0sm_b0m_v0m_n48));
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u138 (.A0(c0sm_b0m_v0m_n350), .A1(c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n166), .C0(c0sm_b0m_v0m_n167), .Y(c0sm_b0m_v0m_n49));
  AOI21_X0P5M_A12TR c0sm_b0m_v0m_u9 (.A0(c0sm_b0m_v0m_n3), .A1(c0nm_b0m_v0m_n4), .B0(c0sm_b0m_v0m_n8), .Y(c0sm_b0m_v0m_n5));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u6 (.A(c0sm_b0m_v0m_n1), .B(c0nm_b0m_v0m_n4), .C(c0sm_b0m_v0m_tail_0_), .Y(c0sm_b0m_v0m_n6));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u223 (.A(c0sm_b0m_v0m_buffers3_7_), .Y(c0sm_b0m_v0m_n62));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u142 (.A(c0sm_b0m_v0m_n169), .Y(c0sm_b0m_v0m_n63));
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u145 (.A0(c0sm_b0m_v0m_n351), .A1(c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n172), .C0(c0sm_b0m_v0m_n173), .Y(c0sm_b0m_v0m_n64));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u218 (.A(c0sm_b0m_v0m_buffers3_8_), .Y(c0sm_b0m_v0m_n65));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u149 (.A(c0sm_b0m_v0m_n175), .Y(c0sm_b0m_v0m_n66));
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u152 (.A0(c0sm_b0m_v0m_n352), .A1(c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n178), .C0(c0sm_b0m_v0m_n179), .Y(c0sm_b0m_v0m_n67));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u213 (.A(c0sm_b0m_v0m_buffers3_9_), .Y(c0sm_b0m_v0m_n68));
  // BSIM@ modules: mx216 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u156 (.A(c0sm_b0m_v0m_n181), .Y(c0sm_b0m_v0m_n69));
  // BSIM@ modules: mx281 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u193 (.A(c0sm_b0m_v0m_tail_1_), .Y(c0sm_b0m_v0m_n7));
  OA211_X0P5M_A12TR c0sm_b0m_v0m_u159 (.A0(c0sm_b0m_v0m_n353), .A1(c0sm_b0m_v0m_n135), .B0(c0sm_b0m_v0m_n184), .C0(c0sm_b0m_v0m_n185), .Y(c0sm_b0m_v0m_n70));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u258 (.A(c0sm_b0m_v0m_buffers3_10_), .Y(c0sm_b0m_v0m_n71));
  // BSIM@ modules: mx281 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u165 (.A(c0sm_b0m_v0m_n26), .Y(c0sm_b0m_v0m_n72));
  AOI21_X0P5M_A12TR c0sm_b0m_v0m_u274 (.A0(c0sm_b0m_v0m_head_0_), .A1(c0sm_b0m_v0m_head_1_), .B0(c0sm_b0m_v0m_head_2_), .Y(c0sm_b0m_v0m_n73));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u36 (.A(c0sm_b0m_v0m_buffers0_0_), .Y(c0sm_b0m_v0m_n74));
  // BSIM@ modules: mx372 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0sm_b0m_v0m_u35 (.A0(c0sm_b0m_v0m_n77), .A1(c0sm_b0m_v0m_n25), .B0(c0sm_b0m_v0m_n78), .B1(c0sm_b0m_v0m_n27), .C0(reset), .Y(c0sm_b0m_v0m_n75));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u62 (.A(c0sm_b0m_v0m_n95), .B(c0nm_b0m_v0m_n4), .C(c0sm_b0m_v0m_n96), .Y(c0sm_b0m_v0m_n76));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u64 (.A(c0sm_b0m_v0m_n95), .Y(c0sm_b0m_v0m_n77));
  // BSIM@ modules: mx281 
  // BSIM@ covered_modules=1 :   NAND3_X0P5A_A12TR c0sm_b0m_v0m_u61 (.A(c0sm_b0m_v0m_n93), .B(c0sm_b0m_v0m_n94), .C(c0sm_b0m_v0m_n72), .Y(c0sm_b0m_v0m_n78));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u39 (.A(c0sm_b0m_v0m_buffers0_1_), .Y(c0sm_b0m_v0m_n79));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0sm_b0m_v0m_u10 (.A(reset), .B(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n8));
  // BSIM@ modules: mx372 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0sm_b0m_v0m_u38 (.A0(c0sm_b0m_v0m_n77), .A1(c0sm_b0m_v0m_n31), .B0(c0sm_b0m_v0m_n78), .B1(c0sm_b0m_v0m_n32), .C0(reset), .Y(c0sm_b0m_v0m_n80));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR c0sm_b0m_v0m_u63 (.A(c0sm_b0m_v0m_n77), .B(c0nm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n81));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u60 (.A(c0sm_b0m_v0m_n76), .B(c0nm_b0m_v0m_n4), .C(c0sm_b0m_v0m_n78), .Y(c0sm_b0m_v0m_n82));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u41 (.A(c0sm_b0m_v0m_buffers0_2_), .Y(c0sm_b0m_v0m_n83));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u43 (.A(c0sm_b0m_v0m_buffers0_3_), .Y(c0sm_b0m_v0m_n84));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u45 (.A(c0sm_b0m_v0m_buffers0_4_), .Y(c0sm_b0m_v0m_n85));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u47 (.A(c0sm_b0m_v0m_buffers0_5_), .Y(c0sm_b0m_v0m_n86));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u49 (.A(c0sm_b0m_v0m_buffers0_6_), .Y(c0sm_b0m_v0m_n87));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u51 (.A(c0sm_b0m_v0m_buffers0_7_), .Y(c0sm_b0m_v0m_n88));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u53 (.A(c0sm_b0m_v0m_buffers0_8_), .Y(c0sm_b0m_v0m_n89));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u55 (.A(c0sm_b0m_v0m_buffers0_9_), .Y(c0sm_b0m_v0m_n90));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u57 (.A(c0sm_b0m_v0m_buffers0_10_), .Y(c0sm_b0m_v0m_n91));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u59 (.A(c0sm_b0m_v0m_buffers0_11_), .Y(c0sm_b0m_v0m_n92));
  // BSIM@ modules: mx281 
  // BSIM@ covered_modules=1 :   NAND3_X0P5A_A12TR c0sm_b0m_v0m_u192 (.A(c0sm_b0m_v0m_tail_0_), .B(c0sm_b0m_v0m_n7), .C(c0sm_b0m_v0m_n355), .Y(c0sm_b0m_v0m_n93));
  // BSIM@ modules: mx281 
  // BSIM@ covered_modules=1 :   NAND3_X0P5A_A12TR c0sm_b0m_v0m_u188 (.A(c0sm_b0m_v0m_tail_1_), .B(c0sm_b0m_v0m_n3), .C(c0sm_b0m_v0m_n355), .Y(c0sm_b0m_v0m_n94));
  // BSIM@ modules: mx281 
  // BSIM@ covered_modules=1 :   NAND3_X0P5A_A12TR c0sm_b0m_v0m_u186 (.A(c0sm_b0m_v0m_n3), .B(c0sm_b0m_v0m_n7), .C(c0sm_b0m_v0m_n355), .Y(c0sm_b0m_v0m_n95));
  // BSIM@ modules: mx316 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u177 (.A(c0sm_b0m_v0m_n193), .Y(c0sm_b0m_v0m_n96));
  // BSIM@ modules: mx132 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0sm_b0m_v0m_u66 (.A0(c0sm_b0m_v0m_n99), .A1(c0sm_b0m_v0m_n25), .B0(c0sm_b0m_v0m_n100), .B1(c0sm_b0m_v0m_n27), .C0(reset), .Y(c0sm_b0m_v0m_n97));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u81 (.A(c0sm_b0m_v0m_n93), .B(c0nm_b0m_v0m_n4), .C(c0sm_b0m_v0m_n104), .Y(c0sm_b0m_v0m_n98));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_b0m_v0m_u83 (.A(c0sm_b0m_v0m_n93), .Y(c0sm_b0m_v0m_n99));
  // BSIM@ modules: mx407 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0sm_b0m_v0m_tail_reg_0_ (.CK(clk), .Q(c0sm_b0m_v0m_tail_0_), .D(c0sm_b0m_v0m_n277));
  // BSIM@ modules: mx407 
  // BSIM@ covered_modules=1 :   DFFQ_X1M_A12TR c0sm_b0m_v0m_tail_reg_1_ (.CK(clk), .Q(c0sm_b0m_v0m_tail_1_), .D(c0sm_b0m_v0m_n278));
  // BSIM@ modules: mx326 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u13 (.A(flitin_1[10]), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_10_));
  // BSIM@ modules: mx326 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u12 (.A(flitin_1[11]), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_11_));
  // BSIM@ modules: mx326 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u11 (.A(flitin_1[2]), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_2_));
  // BSIM@ modules: mx326 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u10 (.A(flitin_1[3]), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_3_));
  // BSIM@ modules: mx326 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u9 (.A(flitin_1[4]), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_4_));
  // BSIM@ modules: mx326 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u8 (.A(flitin_1[5]), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_5_));
  // BSIM@ modules: mx326 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u7 (.A(flitin_1[6]), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_6_));
  // BSIM@ modules: mx326 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u6 (.A(flitin_1[7]), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_7_));
  // BSIM@ modules: mx326 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u5 (.A(flitin_1[8]), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_8_));
  // BSIM@ modules: mx326 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u4 (.A(flitin_1[9]), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_9_));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u268 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n105), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n23), .C0(c0sm_b0m_v0m_n276), .Y(c0sm_headflit[0]));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u263 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n122), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n29), .C0(c0sm_b0m_v0m_n275), .Y(c0sm_headflit[1]));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u245 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n131), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n35), .C0(c0sm_b0m_v0m_n272), .Y(c0sm_headflit[2]));
  // BSIM@ modules: mx212 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u240 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n138), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n38), .C0(c0sm_b0m_v0m_n271), .Y(c0sm_headflit[3]));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u235 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n144), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n41), .C0(c0sm_b0m_v0m_n270), .Y(c0sm_headflit[4]));
  // BSIM@ modules: mx212 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u230 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n150), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n44), .C0(c0sm_b0m_v0m_n269), .Y(c0sm_headflit[5]));
  // BSIM@ modules: mx212 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u225 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n156), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n47), .C0(c0sm_b0m_v0m_n268), .Y(c0sm_headflit[6]));
  // BSIM@ modules: mx387 
  // BSIM@ covered_modules=1 :   OAI221_X0P5M_A12TR c0sm_b0m_v0m_u220 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n162), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n62), .C0(c0sm_b0m_v0m_n267), .Y(c0sm_headflit[7]));
  // BSIM@ modules: mx345 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR c0sm_u3 (.A(flitin_1[1]), .B(flitin_1[0]), .Y(c0sm_n3));
  NOR2B_X0P5M_A12TR c0sm_u4 (.AN(c0sm_headflit[1]), .B(c0sm_headflit[0]), .Y(c0sm_n4));
  INV_X0P5B_A12TR c0sm_r0m_u6 (.A(c0sm_n4), .Y(c0sm_r0m_n1));
  AOI2XB1_X0P5M_A12TR c0sm_r0m_u10 (.A0(curry[2]), .A1N(c0sm_headflit[4]), .B0(c0sm_r0m_n11), .Y(c0sm_r0m_n10));
  NOR3_X0P5A_A12TR c0sm_r0m_u5 (.A(c0sm_r0m_n3), .B(reset), .C(c0sm_r0m_n1), .Y(c0sm_r0m_n100));
  AOI2XB1_X0P5M_A12TR c0sm_r0m_u11 (.A0(c0sm_headflit[4]), .A1N(curry[2]), .B0(c0sm_r0m_n12), .Y(c0sm_r0m_n11));
  NOR3_X0P5A_A12TR c0sm_r0m_u3 (.A(c0sm_r0m_n1), .B(reset), .C(c0sm_r0m_n2), .Y(c0sm_r0m_n110));
  // BSIM@ modules: mx29 
  // BSIM@ covered_modules=1 :   AOI22_X0P5M_A12TR c0sm_r0m_u12 (.A0(c0sm_r0m_n13), .A1(curry[0]), .B0(curry[1]), .B1(c0sm_r0m_n14), .Y(c0sm_r0m_n12));
  AOI2XB1_X0P5M_A12TR c0sm_r0m_u14 (.A0(c0sm_headflit[3]), .A1N(curry[1]), .B0(c0sm_headflit[2]), .Y(c0sm_r0m_n13));
  // BSIM@ modules: mx212 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_r0m_u13 (.A(c0sm_headflit[3]), .Y(c0sm_r0m_n14));
  // BSIM@ modules: mx334 
  // BSIM@ covered_modules=1 :   OR2_X0P5M_A12TR c0sm_r0m_u18 (.A(currx[0]), .B(c0sm_r0m_n9), .Y(c0sm_r0m_n15));
  // BSIM@ modules: mx319 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_r0m_u16 (.A(c0sm_r0m_n15), .B(currx[1]), .Y(c0sm_r0m_n16));
  INV_X0P5B_A12TR c0sm_r0m_u4 (.A(c0sm_r0m_n3), .Y(c0sm_r0m_n2));
  AO1B2_X0P5M_A12TR c0sm_r0m_u7 (.A0N(c0sm_r0m_n5), .B0(c0nm_r0m_n4), .B1(c0sm_headflit[7]), .Y(c0sm_r0m_n3));
  OAI22_X0P5M_A12TR c0sm_r0m_u8 (.A0(c0sm_r0m_n6), .A1(c0sm_r0m_n7), .B0(c0sm_headflit[7]), .B1(c0nm_r0m_n4), .Y(c0sm_r0m_n5));
  OA21A1OI2_X0P5M_A12TR c0sm_r0m_u15 (.A0(currx[1]), .A1(c0sm_r0m_n15), .B0(c0sm_r0m_n8), .C0(c0sm_r0m_n16), .Y(c0sm_r0m_n6));
  // BSIM@ modules: mx110 
  // BSIM@ covered_modules=1 :   AOI221_X0P5M_A12TR c0sm_r0m_u9 (.A0(currx[1]), .A1(c0sm_r0m_n8), .B0(currx[0]), .B1(c0sm_r0m_n9), .C0(c0sm_r0m_n10), .Y(c0sm_r0m_n7));
  // BSIM@ modules: mx212 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_r0m_u17 (.A(c0sm_headflit[6]), .Y(c0sm_r0m_n8));
  // BSIM@ modules: mx212 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_r0m_u19 (.A(c0sm_headflit[5]), .Y(c0sm_r0m_n9));
  DFFQ_X1M_A12TR c0sm_r0m_vc_req_reg_0_ (.CK(clk), .Q(c0sm_routewire[0]), .D(c0sm_r0m_n100));
  DFFQ_X1M_A12TR c0sm_r0m_vc_req_reg_1_ (.CK(clk), .Q(c0sm_routewire[1]), .D(c0sm_r0m_n110));
  DFFQ_X1M_A12TR c0sm_v0m_full_reg (.CK(clk), .Q(c0sm_v0m_full), .D(c0sm_v0m_n64));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_v0m_u9 (.A(c0sm_v0m_n8), .Y(c0sm_v0m_n1));
  AOI32_X0P5M_A12TR c0sm_v0m_u12 (.A0(c0sm_v0m_n11), .A1(c0sm_v0m_n9), .A2(c0sm_n3), .B0(c0sm_v0m_full), .B1(c0sm_v0m_n12), .Y(c0sm_v0m_n10));
  INV_X0P5B_A12TR c0sm_v0m_u14 (.A(c0sm_v0m_n14), .Y(c0sm_v0m_n11));
  INV_X0P5B_A12TR c0sm_v0m_u13 (.A(c0sm_v0m_n13), .Y(c0sm_v0m_n12));
  // BSIM@ modules: mx361 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0sm_v0m_u30 (.A(c0sm_v0m_n9), .B(c0sm_n3), .Y(c0sm_v0m_n13));
  NAND3_X0P5A_A12TR c0sm_v0m_u28 (.A(c0sm_v0m_state_queuelen_0_), .B(c0sm_v0m_n17), .C(c0sm_v0m_state_queuelen_1_), .Y(c0sm_v0m_n14));
  // BSIM@ modules: mx22 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0sm_v0m_u16 (.A(c0sm_v0m_state_queuelen_0_), .B(c0sm_v0m_n18), .S0(c0sm_v0m_state_queuelen_1_), .Y(c0sm_v0m_n15));
  AOI21_X0P5M_A12TR c0sm_v0m_u20 (.A0(c0sm_v0m_n23), .A1(c0sm_v0m_n22), .B0(c0sm_v0m_n24), .Y(c0sm_v0m_n16));
  INV_X0P5B_A12TR c0sm_v0m_u29 (.A(c0sm_v0m_state_queuelen_2_), .Y(c0sm_v0m_n17));
  NAND3_X0P5A_A12TR c0sm_v0m_u27 (.A(c0sm_v0m_n14), .B(c0sm_v0m_n9), .C(c0sm_n3), .Y(c0sm_v0m_n18));
  // BSIM@ modules: mx22 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0sm_v0m_u18 (.A(c0sm_v0m_n20), .B(c0sm_v0m_n21), .S0(c0sm_v0m_state_queuelen_1_), .Y(c0sm_v0m_n19));
  // BSIM@ modules: mx21 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0sm_v0m_u4 (.A(c0sm_v0m_n3), .B(c0sm_routewire[1]), .S0(c0sm_v0m_n4), .Y(c0sm_v0m_n2));
  MXIT2_X0P5M_A12TR c0sm_v0m_u21 (.A(c0sm_v0m_n18), .B(c0sm_v0m_n25), .S0(c0sm_v0m_n23), .Y(c0sm_v0m_n20));
  OAI21_X0P5M_A12TR c0sm_v0m_u19 (.A0(c0sm_v0m_n22), .A1(c0sm_v0m_n23), .B0(c0sm_v0m_n16), .Y(c0sm_v0m_n21));
  INV_X0P5B_A12TR c0sm_v0m_u26 (.A(c0sm_v0m_n18), .Y(c0sm_v0m_n22));
  INV_X0P5B_A12TR c0sm_v0m_u34 (.A(c0sm_v0m_state_queuelen_0_), .Y(c0sm_v0m_n23));
  AOI21_X0P5M_A12TR c0sm_v0m_u25 (.A0(c0sm_v0m_n26), .A1(c0sm_v0m_n13), .B0(c0sm_v0m_n22), .Y(c0sm_v0m_n24));
  NAND2_X0P5A_A12TR c0sm_v0m_u22 (.A(c0sm_v0m_n13), .B(c0sm_v0m_n26), .Y(c0sm_v0m_n25));
  INV_X0P5B_A12TR c0sm_v0m_u33 (.A(c0sm_v0m_full), .Y(c0sm_v0m_n26));
  XNOR2_X0P5M_A12TR c0sm_v0m_u24 (.A(c0sm_v0m_n23), .B(c0sm_v0m_n24), .Y(c0sm_v0m_n27));
  OAI31_X0P5M_A12TR c0sm_v0m_u32 (.A0(c0sm_v0m_n29), .A1(tailout_1), .A2(c0sm_v0m_state_status_0_), .B0(c0sm_v0m_n5), .Y(c0sm_v0m_n28));
  INV_X0P5B_A12TR c0sm_v0m_u40 (.A(c0sm_v0m_state_status_1_), .Y(c0sm_v0m_n29));
  // BSIM@ modules: mx330 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_v0m_u5 (.A(swalloc_req_1[1]), .B(c0sm_v0m_n5), .Y(c0sm_v0m_n3));
  // BSIM@ modules: mx363 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0sm_v0m_u3 (.A(c0sm_v0m_n1), .B(c0sm_v0m_n2), .Y(c0sm_v0m_n32));
  // BSIM@ modules: mx363 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0sm_v0m_u6 (.A(c0sm_v0m_n1), .B(c0sm_v0m_n6), .Y(c0sm_v0m_n33));
  OA211_X0P5M_A12TR c0sm_v0m_u36 (.A0(c0sm_routewire[1]), .A1(c0sm_routewire[0]), .B0(c0sm_v0m_state_status_0_), .C0(c0sm_v0m_state_status_1_), .Y(c0sm_v0m_n4));
  OAI211_X0P5M_A12TR c0sm_v0m_u39 (.A0(swalloc_resp_1[1]), .A1(swalloc_resp_1[0]), .B0(c0sm_v0m_n29), .C0(c0sm_v0m_state_status_0_), .Y(c0sm_v0m_n5));
  AO1B2_X0P5M_A12TR c0sm_v0m_u37 (.A0N(c0sm_v0m_n8), .B0(c0sm_v0m_n5), .B1(c0sm_v0m_state_status_0_), .Y(c0sm_v0m_n57));
  AO21A1AI2_X0P5M_A12TR c0sm_v0m_u35 (.A0(c0sm_v0m_n29), .A1(c0sm_v0m_n5), .B0(c0sm_v0m_n4), .C0(c0sm_v0m_n8), .Y(c0sm_v0m_n58));
  // BSIM@ modules: mx21 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR c0sm_v0m_u7 (.A(c0sm_v0m_n7), .B(c0sm_routewire[0]), .S0(c0sm_v0m_n4), .Y(c0sm_v0m_n6));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0sm_v0m_u23 (.A(reset), .B(c0sm_v0m_n27), .Y(c0sm_v0m_n61));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0sm_v0m_u17 (.A(reset), .B(c0sm_v0m_n19), .Y(c0sm_v0m_n62));
  AOI211_X0P5M_A12TR c0sm_v0m_u15 (.A0(c0sm_v0m_n15), .A1(c0sm_v0m_n16), .B0(c0sm_v0m_n17), .C0(reset), .Y(c0sm_v0m_n63));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0sm_v0m_u11 (.A(reset), .B(c0sm_v0m_n10), .Y(c0sm_v0m_n64));
  // BSIM@ modules: mx331 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_v0m_u8 (.A(swalloc_req_1[0]), .B(c0sm_v0m_n5), .Y(c0sm_v0m_n7));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR c0sm_v0m_u38 (.A(reset), .B(tailout_1), .Y(c0sm_v0m_n8));
  OAI31_X0P5M_A12TR c0sm_v0m_u31 (.A0(c0sm_v0m_state_queuelen_0_), .A1(c0sm_v0m_state_queuelen_2_), .A2(c0sm_v0m_state_queuelen_1_), .B0(c0sm_v0m_n28), .Y(c0sm_v0m_n9));
  DFFQ_X1M_A12TR c0sm_v0m_state_queuelen_reg_0_ (.CK(clk), .Q(c0sm_v0m_state_queuelen_0_), .D(c0sm_v0m_n61));
  DFFQ_X1M_A12TR c0sm_v0m_state_queuelen_reg_1_ (.CK(clk), .Q(c0sm_v0m_state_queuelen_1_), .D(c0sm_v0m_n62));
  DFFQ_X1M_A12TR c0sm_v0m_state_queuelen_reg_2_ (.CK(clk), .Q(c0sm_v0m_state_queuelen_2_), .D(c0sm_v0m_n63));
  DFFQ_X1M_A12TR c0sm_v0m_state_status_reg_0_ (.CK(clk), .Q(c0sm_v0m_state_status_0_), .D(c0sm_v0m_n57));
  DFFQ_X1M_A12TR c0sm_v0m_state_status_reg_1_ (.CK(clk), .Q(c0sm_v0m_state_status_1_), .D(c0sm_v0m_n58));
  // BSIM@ modules: mx259 
  // BSIM@ covered_modules=1 :   NAND2B_X0P5M_A12TR d0m_u2 (.AN(swalloc_resp_1[0]), .B(swalloc_resp_0[0]), .Y(colsel0[0]));
  // BSIM@ modules: mx259 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR d0m_u1 (.A(swalloc_resp_1[0]), .B(swalloc_resp_0[0]), .Y(colsel0[1]));
  // BSIM@ modules: mx260 
  // BSIM@ covered_modules=1 :   NAND2B_X0P5M_A12TR d1m_u2 (.AN(swalloc_resp_1[1]), .B(swalloc_resp_0[1]), .Y(colsel1[0]));
  // BSIM@ modules: mx260 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR d1m_u1 (.A(swalloc_resp_1[1]), .B(swalloc_resp_0[1]), .Y(colsel1[1]));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2B_X0P5M_A12TR c0nm_u5 (.AN(debitout_0), .B(reset), .Y(creditout_0));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2B_X0P5M_A12TR c0sm_u5 (.AN(debitout_1), .B(reset), .Y(creditout_1));
  // BSIM@ modules: mx356 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0nm_v0m_u10 (.A(c0nm_v0m_n9), .Y(debitout_0));
  // BSIM@ modules: mx361 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR c0sm_v0m_u10 (.A(c0sm_v0m_n9), .Y(debitout_1));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx0m_m0m_m4m_u1 (.A(x0m_bx0m_m0m_int01), .B(x0m__logic1_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[0]));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx10m_m0m_m4m_u1 (.A(x0m_bx10m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[10]));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx11m_m0m_m4m_u1 (.A(x0m_bx11m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[11]));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx1m_m0m_m4m_u1 (.A(x0m_bx1m_m0m_int01), .B(x0m__logic1_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[1]));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx2m_m0m_m4m_u1 (.A(x0m_bx2m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[2]));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx3m_m0m_m4m_u1 (.A(x0m_bx3m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[3]));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx4m_m0m_m4m_u1 (.A(x0m_bx4m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[4]));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx5m_m0m_m4m_u1 (.A(x0m_bx5m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[5]));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx6m_m0m_m4m_u1 (.A(x0m_bx6m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[6]));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx7m_m0m_m4m_u1 (.A(x0m_bx7m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[7]));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx8m_m0m_m4m_u1 (.A(x0m_bx8m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[8]));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx9m_m0m_m4m_u1 (.A(x0m_bx9m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0[9]));
  // BSIM@ modules: mx341 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx0m_m1m_m4m_u1 (.A(x0m_bx0m_m1m_int01), .B(x0m__logic1_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[0]));
  // BSIM@ modules: mx101 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx10m_m1m_m4m_u1 (.A(x0m_bx10m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[10]));
  // BSIM@ modules: mx10 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx11m_m1m_m4m_u1 (.A(x0m_bx11m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[11]));
  // BSIM@ modules: mx341 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx1m_m1m_m4m_u1 (.A(x0m_bx1m_m1m_int01), .B(x0m__logic1_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[1]));
  // BSIM@ modules: mx101 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx2m_m1m_m4m_u1 (.A(x0m_bx2m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[2]));
  // BSIM@ modules: mx101 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx3m_m1m_m4m_u1 (.A(x0m_bx3m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[3]));
  // BSIM@ modules: mx10 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx4m_m1m_m4m_u1 (.A(x0m_bx4m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[4]));
  // BSIM@ modules: mx101 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx5m_m1m_m4m_u1 (.A(x0m_bx5m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[5]));
  // BSIM@ modules: mx101 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx6m_m1m_m4m_u1 (.A(x0m_bx6m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[6]));
  // BSIM@ modules: mx101 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx7m_m1m_m4m_u1 (.A(x0m_bx7m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[7]));
  // BSIM@ modules: mx101 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx8m_m1m_m4m_u1 (.A(x0m_bx8m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[8]));
  // BSIM@ modules: mx101 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx9m_m1m_m4m_u1 (.A(x0m_bx9m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1[9]));
  NAND2B_X0P5M_A12TR c0nm_b0m_u26 (.AN(c0nm_b0m_rdata[0]), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0[0]));
  // BSIM@ modules: mx321 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u25 (.A(c0nm_b0m_rdata[10]), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0[10]));
  // BSIM@ modules: mx321 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u24 (.A(c0nm_b0m_rdata[11]), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0[11]));
  NAND2B_X0P5M_A12TR c0nm_b0m_u23 (.AN(c0nm_b0m_rdata[1]), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0[1]));
  // BSIM@ modules: mx321 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u22 (.A(c0nm_b0m_rdata[2]), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0[2]));
  // BSIM@ modules: mx321 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u21 (.A(c0nm_b0m_rdata[3]), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0[3]));
  // BSIM@ modules: mx321 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u20 (.A(c0nm_b0m_rdata[4]), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0[4]));
  // BSIM@ modules: mx321 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u19 (.A(c0nm_b0m_rdata[5]), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0[5]));
  // BSIM@ modules: mx321 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u18 (.A(c0nm_b0m_rdata[6]), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0[6]));
  // BSIM@ modules: mx321 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u17 (.A(c0nm_b0m_rdata[7]), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0[7]));
  // BSIM@ modules: mx321 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u16 (.A(c0nm_b0m_rdata[8]), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0[8]));
  // BSIM@ modules: mx321 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0nm_b0m_u15 (.A(c0nm_b0m_rdata[9]), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0[9]));
  NAND2B_X0P5M_A12TR c0sm_b0m_u26 (.AN(c0sm_b0m_rdata[0]), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1[0]));
  // BSIM@ modules: mx327 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u25 (.A(c0sm_b0m_rdata[10]), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1[10]));
  // BSIM@ modules: mx327 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u24 (.A(c0sm_b0m_rdata[11]), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1[11]));
  NAND2B_X0P5M_A12TR c0sm_b0m_u23 (.AN(c0sm_b0m_rdata[1]), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1[1]));
  // BSIM@ modules: mx327 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u22 (.A(c0sm_b0m_rdata[2]), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1[2]));
  // BSIM@ modules: mx327 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u21 (.A(c0sm_b0m_rdata[3]), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1[3]));
  // BSIM@ modules: mx327 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u20 (.A(c0sm_b0m_rdata[4]), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1[4]));
  // BSIM@ modules: mx327 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u19 (.A(c0sm_b0m_rdata[5]), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1[5]));
  // BSIM@ modules: mx327 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u18 (.A(c0sm_b0m_rdata[6]), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1[6]));
  // BSIM@ modules: mx327 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u17 (.A(c0sm_b0m_rdata[7]), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1[7]));
  // BSIM@ modules: mx327 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u16 (.A(c0sm_b0m_rdata[8]), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1[8]));
  // BSIM@ modules: mx327 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR c0sm_b0m_u15 (.A(c0sm_b0m_rdata[9]), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1[9]));
  TIELO_X1M_A12TR u1 (.Y(net1));
  // BSIM@ modules: mx25 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR s0m_u13 (.A(s0m_n4), .B(s0m_n5), .S0(s0m_state_invc0_0_), .Y(nomorebufs_0));
  MXIT2_X0P5M_A12TR s0m_u12 (.A(s0m_n4), .B(s0m_n5), .S0(s0m_state_invc0_1_), .Y(nomorebufs_1));
  // BSIM@ modules: mx5 
  // BSIM@ covered_modules=1 :   TIELO_X1M_A12TR s0m_u2 (.Y(s0m__logic0_));
  // BSIM@ modules: mx25 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR s0m_u36 (.A(s0m_n26), .B(c0nm_v0m_n9), .S0(s0m_state_invc0_0_), .Y(s0m_debit_outvc0));
  // BSIM@ modules: mx26 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR s0m_u34 (.A(s0m_n20), .B(c0nm_v0m_n9), .S0(s0m_state_invc1_0_), .Y(s0m_debit_outvc1));
  DFFQ_X1M_A12TR s0m_o0nm_eligible_reg (.CK(clk), .Q(s0m_elig_0_), .D(s0m_o0nm_n41));
  DFFQ_X1M_A12TR s0m_o0sm_eligible_reg (.CK(clk), .Q(s0m_elig_1_), .D(s0m_o0sm_n41));
  INV_X0P5B_A12TR s0m_m0m_u8 (.A(s0m_request0[0]), .Y(s0m_m0m_n1));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR s0m_m0m_u4 (.A(reset), .B(s0m_m0m_n2), .Y(s0m_m0m_n10));
  // BSIM@ modules: mx5 
  // BSIM@ covered_modules=1 :   XOR2_X0P5M_A12TR s0m_m0m_u5 (.A(s0m__logic0_), .B(s0m_m0m_n3), .Y(s0m_m0m_n2));
  // BSIM@ modules: mx5 
  // BSIM@ covered_modules=1 :   AOI2XB1_X0P5M_A12TR s0m_m0m_u6 (.A0(s0m_m0m_row1_0_), .A1N(s0m_request1[0]), .B0(s0m_outb0_0_), .Y(s0m_m0m_n3));
  DFFQ_X1M_A12TR s0m_m0m_state1_reg (.CK(clk), .Q(s0m_m0m_row1_0_), .D(s0m_m0m_n10));
  INV_X0P5B_A12TR s0m_m1m_u8 (.A(s0m_request0[1]), .Y(s0m_m1m_n1));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR s0m_m1m_u4 (.A(reset), .B(s0m_m1m_n2), .Y(s0m_m1m_n10));
  XOR2_X0P5M_A12TR s0m_m1m_u5 (.A(s0m__logic0_), .B(s0m_m1m_n3), .Y(s0m_m1m_n2));
  AOI2XB1_X0P5M_A12TR s0m_m1m_u6 (.A0(s0m_m1m_row1_0_), .A1N(s0m_request1[1]), .B0(s0m_outb1_0_), .Y(s0m_m1m_n3));
  DFFQ_X1M_A12TR s0m_m1m_state1_reg (.CK(clk), .Q(s0m_m1m_row1_0_), .D(s0m_m1m_n10));
  // BSIM@ modules: mx347 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR s0m_u4 (.A(tailout_1), .B(s0m_state_invc1_1_), .Y(s0m_n1));
  INV_X0P5B_A12TR s0m_u24 (.A(swalloc_resp_0[1]), .Y(s0m_n10));
  // BSIM@ modules: mx350 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR s0m_u22 (.A(s0m_outb1_0_), .B(s0m_n9), .Y(s0m_n11));
  NOR2_X0P5A_A12TR s0m_u21 (.A(swalloc_req_0[1]), .B(swalloc_req_0[0]), .Y(s0m_n12));
  INV_X0P5B_A12TR s0m_u27 (.A(swalloc_resp_1[0]), .Y(s0m_n13));
  // BSIM@ modules: mx349 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR s0m_u26 (.A(s0m_outb0_1_), .B(s0m_n16), .Y(s0m_n14));
  OAI31_X0P5M_A12TR s0m_u29 (.A0(s0m_n19), .A1(swalloc_resp_1[1]), .A2(swalloc_resp_1[0]), .B0(s0m_n16), .Y(s0m_n15));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR s0m_u32 (.A(reset), .B(tailout_1), .Y(s0m_n16));
  INV_X0P5B_A12TR s0m_u33 (.A(swalloc_resp_1[1]), .Y(s0m_n17));
  // BSIM@ modules: mx349 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR s0m_u31 (.A(s0m_outb1_1_), .B(s0m_n16), .Y(s0m_n18));
  NOR2_X0P5A_A12TR s0m_u30 (.A(swalloc_req_1[1]), .B(swalloc_req_1[0]), .Y(s0m_n19));
  INV_X0P5B_A12TR s0m_u6 (.A(tailout_0), .Y(s0m_n2));
  // BSIM@ modules: mx348 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR s0m_u35 (.A(debitout_1), .B(s0m_state_invc1_1_), .Y(s0m_n20));
  // BSIM@ modules: mx23 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR s0m_u28 (.A(s0m_n17), .B(s0m_n18), .S0(s0m_n15), .Y(s0m_n22));
  // BSIM@ modules: mx23 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR s0m_u25 (.A(s0m_n13), .B(s0m_n14), .S0(s0m_n15), .Y(s0m_n23));
  // BSIM@ modules: mx24 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR s0m_u19 (.A(s0m_n10), .B(s0m_n11), .S0(s0m_n8), .Y(s0m_n24));
  // BSIM@ modules: mx24 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR s0m_u16 (.A(s0m_n6), .B(s0m_n7), .S0(s0m_n8), .Y(s0m_n25));
  // BSIM@ modules: mx348 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR s0m_u38 (.A(debitout_1), .B(s0m_state_invc0_1_), .Y(s0m_n26));
  // BSIM@ modules: mx347 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR s0m_u7 (.A(s0m_state_invc0_1_), .B(tailout_1), .Y(s0m_n3));
  INV_X0P5B_A12TR s0m_u15 (.A(s0m_no_bufs1), .Y(s0m_n4));
  INV_X0P5B_A12TR s0m_u14 (.A(s0m_no_bufs0), .Y(s0m_n5));
  INV_X0P5B_A12TR s0m_u18 (.A(swalloc_resp_0[0]), .Y(s0m_n6));
  // BSIM@ modules: mx350 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR s0m_u17 (.A(s0m_outb0_0_), .B(s0m_n9), .Y(s0m_n7));
  OAI31_X0P5M_A12TR s0m_u20 (.A0(s0m_n12), .A1(swalloc_resp_0[1]), .A2(swalloc_resp_0[0]), .B0(s0m_n9), .Y(s0m_n8));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR s0m_u23 (.A(reset), .B(tailout_0), .Y(s0m_n9));
  DFFQ_X1M_A12TR s0m_o0nm_no_bufs_reg (.CK(clk), .Q(s0m_no_bufs0), .D(s0m_o0nm_n42));
  DFFQ_X1M_A12TR s0m_o0sm_no_bufs_reg (.CK(clk), .Q(s0m_no_bufs1), .D(s0m_o0sm_n42));
  AO21A1AI2_X0P5M_A12TR s0m_o0nm_u4 (.A0(s0m_o0nm_n2), .A1(s0m_state_invc0_1_), .B0(s0m_outb0_1_), .C0(s0m_o0nm_n3), .Y(s0m_o0nm_n1));
  // BSIM@ modules: mx271 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR s0m_o0nm_u13 (.A(s0m_o0nm_n12), .Y(s0m_o0nm_n11));
  NOR2_X0P5A_A12TR s0m_o0nm_u28 (.A(s0m_o0nm_state_credits_2_), .B(s0m_o0nm_n22), .Y(s0m_o0nm_n12));
  MXIT2_X0P5M_A12TR s0m_o0nm_u15 (.A(s0m_o0nm_n14), .B(s0m_o0nm_n15), .S0(s0m_o0nm_state_credits_2_), .Y(s0m_o0nm_n13));
  NOR3_X0P5A_A12TR s0m_o0nm_u18 (.A(s0m_o0nm_n18), .B(s0m_o0nm_n20), .C(s0m_o0nm_n16), .Y(s0m_o0nm_n14));
  NAND2B_X0P5M_A12TR s0m_o0nm_u16 (.AN(s0m_o0nm_n16), .B(s0m_o0nm_n17), .Y(s0m_o0nm_n15));
  NOR2_X0P5A_A12TR s0m_o0nm_u26 (.A(s0m_o0nm_n23), .B(s0m_o0nm_n20), .Y(s0m_o0nm_n16));
  XOR2_X0P5M_A12TR s0m_o0nm_u17 (.A(s0m_o0nm_n18), .B(s0m_o0nm_n19), .Y(s0m_o0nm_n17));
  // BSIM@ modules: mx261 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR s0m_o0nm_u22 (.A(s0m_o0nm_state_credits_1_), .B(s0m_o0nm_state_credits_0_), .Y(s0m_o0nm_n18));
  AO1B2_X0P5M_A12TR s0m_o0nm_u21 (.A0N(s0m_o0nm_n20), .B0(s0m_o0nm_n18), .B1(s0m_o0nm_n22), .Y(s0m_o0nm_n19));
  INV_X0P5B_A12TR s0m_o0nm_u5 (.A(s0m_outb0_0_), .Y(s0m_o0nm_n2));
  // BSIM@ modules: mx271 
  // BSIM@ covered_modules=1 :   NOR3_X0P5A_A12TR s0m_o0nm_u27 (.A(s0m_o0nm_n9), .B(creditin_0), .C(s0m_o0nm_n12), .Y(s0m_o0nm_n20));
  AOI32_X0P5M_A12TR s0m_o0nm_u20 (.A0(s0m_o0nm_n22), .A1(s0m_o0nm_n18), .A2(s0m_o0nm_n23), .B0(s0m_o0nm_n16), .B1(s0m_o0nm_state_credits_1_), .Y(s0m_o0nm_n21));
  // BSIM@ modules: mx261 
  // BSIM@ covered_modules=1 :   OR2_X0P5M_A12TR s0m_o0nm_u29 (.A(s0m_o0nm_state_credits_1_), .B(s0m_o0nm_state_credits_0_), .Y(s0m_o0nm_n22));
  AND3_X0P5M_A12TR s0m_o0nm_u30 (.A(s0m_o0nm_n9), .B(s0m_n5), .C(creditin_0), .Y(s0m_o0nm_n23));
  XOR2_X0P5M_A12TR s0m_o0nm_u25 (.A(s0m_o0nm_state_credits_0_), .B(s0m_o0nm_n16), .Y(s0m_o0nm_n24));
  OAI31_X0P5M_A12TR s0m_o0nm_u34 (.A0(s0m_outb0_0_), .A1(s0m_o0nm_state_assigned), .A2(s0m_outb0_1_), .B0(s0m_o0nm_n3), .Y(s0m_o0nm_n25));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR s0m_o0nm_u35 (.A(s0m_tail_outvc0), .B(reset), .Y(s0m_o0nm_n3));
  INV_X0P5B_A12TR s0m_o0nm_u6 (.A(s0m_o0nm_n4), .Y(s0m_o0nm_n30));
  INV_X0P5B_A12TR s0m_o0nm_u3 (.A(s0m_o0nm_n1), .Y(s0m_o0nm_n31));
  INV_X0P5B_A12TR s0m_o0nm_u33 (.A(s0m_o0nm_n25), .Y(s0m_o0nm_n35));
  // BSIM@ modules: mx346 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR s0m_o0nm_u23 (.A(s0m_o0nm_n24), .B(c0nm_b0m_v0m_n4), .Y(s0m_o0nm_n36));
  NAND3_X0P5A_A12TR s0m_o0nm_u19 (.A(s0m_o0nm_n19), .B(c0nm_b0m_v0m_n4), .C(s0m_o0nm_n21), .Y(s0m_o0nm_n37));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR s0m_o0nm_u14 (.A(reset), .B(s0m_o0nm_n13), .Y(s0m_o0nm_n38));
  AO21A1AI2_X0P5M_A12TR s0m_o0nm_u7 (.A0(s0m_o0nm_n5), .A1(s0m_state_invc0_0_), .B0(s0m_outb0_0_), .C0(s0m_o0nm_n3), .Y(s0m_o0nm_n4));
  NOR2_X0P5A_A12TR s0m_o0nm_u9 (.A(s0m_o0nm_n42), .B(s0m_o0nm_n35), .Y(s0m_o0nm_n41));
  OA21_X0P5M_A12TR s0m_o0nm_u10 (.A0(s0m_o0nm_n6), .A1(s0m_o0nm_n7), .B0(c0nm_b0m_v0m_n4), .Y(s0m_o0nm_n42));
  INV_X0P5B_A12TR s0m_o0nm_u8 (.A(s0m_outb0_1_), .Y(s0m_o0nm_n5));
  // BSIM@ modules: mx271 
  // BSIM@ covered_modules=1 :   NOR3_X0P5A_A12TR s0m_o0nm_u12 (.A(s0m_o0nm_n11), .B(creditin_0), .C(s0m_o0nm_n9), .Y(s0m_o0nm_n6));
  AOI21_X0P5M_A12TR s0m_o0nm_u11 (.A0(creditin_0), .A1(s0m_o0nm_n9), .B0(s0m_n5), .Y(s0m_o0nm_n7));
  NOR3_X0P5A_A12TR s0m_o0nm_u32 (.A(s0m_outb0_1_), .B(s0m_outb0_0_), .C(s0m_debit_outvc0), .Y(s0m_o0nm_n9));
  DFFQ_X1M_A12TR s0m_o0nm_state_assigned_reg (.CK(clk), .Q(s0m_o0nm_state_assigned), .D(s0m_o0nm_n35));
  DFFQ_X1M_A12TR s0m_o0nm_state_credits_reg_0_ (.CK(clk), .Q(s0m_o0nm_state_credits_0_), .D(s0m_o0nm_n36));
  DFFQ_X1M_A12TR s0m_o0nm_state_credits_reg_1_ (.CK(clk), .Q(s0m_o0nm_state_credits_1_), .D(s0m_o0nm_n37));
  DFFQ_X1M_A12TR s0m_o0nm_state_credits_reg_2_ (.CK(clk), .Q(s0m_o0nm_state_credits_2_), .D(s0m_o0nm_n38));
  AO21A1AI2_X0P5M_A12TR s0m_o0sm_u4 (.A0(s0m_o0sm_n2), .A1(s0m_state_invc1_1_), .B0(s0m_outb1_1_), .C0(s0m_o0sm_n3), .Y(s0m_o0sm_n1));
  // BSIM@ modules: mx272 
  // BSIM@ covered_modules=1 :   INV_X0P5B_A12TR s0m_o0sm_u13 (.A(s0m_o0sm_n12), .Y(s0m_o0sm_n11));
  NOR2_X0P5A_A12TR s0m_o0sm_u28 (.A(s0m_o0sm_state_credits_2_), .B(s0m_o0sm_n22), .Y(s0m_o0sm_n12));
  MXIT2_X0P5M_A12TR s0m_o0sm_u15 (.A(s0m_o0sm_n14), .B(s0m_o0sm_n15), .S0(s0m_o0sm_state_credits_2_), .Y(s0m_o0sm_n13));
  NOR3_X0P5A_A12TR s0m_o0sm_u18 (.A(s0m_o0sm_n18), .B(s0m_o0sm_n20), .C(s0m_o0sm_n16), .Y(s0m_o0sm_n14));
  NAND2B_X0P5M_A12TR s0m_o0sm_u16 (.AN(s0m_o0sm_n16), .B(s0m_o0sm_n17), .Y(s0m_o0sm_n15));
  NOR2_X0P5A_A12TR s0m_o0sm_u26 (.A(s0m_o0sm_n23), .B(s0m_o0sm_n20), .Y(s0m_o0sm_n16));
  XOR2_X0P5M_A12TR s0m_o0sm_u17 (.A(s0m_o0sm_n18), .B(s0m_o0sm_n19), .Y(s0m_o0sm_n17));
  // BSIM@ modules: mx262 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR s0m_o0sm_u22 (.A(s0m_o0sm_state_credits_1_), .B(s0m_o0sm_state_credits_0_), .Y(s0m_o0sm_n18));
  AO1B2_X0P5M_A12TR s0m_o0sm_u21 (.A0N(s0m_o0sm_n20), .B0(s0m_o0sm_n18), .B1(s0m_o0sm_n22), .Y(s0m_o0sm_n19));
  INV_X0P5B_A12TR s0m_o0sm_u5 (.A(s0m_outb1_0_), .Y(s0m_o0sm_n2));
  // BSIM@ modules: mx272 
  // BSIM@ covered_modules=1 :   NOR3_X0P5A_A12TR s0m_o0sm_u27 (.A(s0m_o0sm_n9), .B(creditin_1), .C(s0m_o0sm_n12), .Y(s0m_o0sm_n20));
  AOI32_X0P5M_A12TR s0m_o0sm_u20 (.A0(s0m_o0sm_n22), .A1(s0m_o0sm_n18), .A2(s0m_o0sm_n23), .B0(s0m_o0sm_n16), .B1(s0m_o0sm_state_credits_1_), .Y(s0m_o0sm_n21));
  // BSIM@ modules: mx262 
  // BSIM@ covered_modules=1 :   OR2_X0P5M_A12TR s0m_o0sm_u29 (.A(s0m_o0sm_state_credits_1_), .B(s0m_o0sm_state_credits_0_), .Y(s0m_o0sm_n22));
  AND3_X0P5M_A12TR s0m_o0sm_u30 (.A(s0m_o0sm_n9), .B(s0m_n4), .C(creditin_1), .Y(s0m_o0sm_n23));
  XOR2_X0P5M_A12TR s0m_o0sm_u25 (.A(s0m_o0sm_state_credits_0_), .B(s0m_o0sm_n16), .Y(s0m_o0sm_n24));
  OAI31_X0P5M_A12TR s0m_o0sm_u34 (.A0(s0m_outb1_0_), .A1(s0m_o0sm_state_assigned), .A2(s0m_outb1_1_), .B0(s0m_o0sm_n3), .Y(s0m_o0sm_n25));
  INV_X0P5B_A12TR s0m_o0sm_u3 (.A(s0m_o0sm_n1), .Y(s0m_o0sm_n26));
  INV_X0P5B_A12TR s0m_o0sm_u6 (.A(s0m_o0sm_n4), .Y(s0m_o0sm_n27));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR s0m_o0sm_u35 (.A(s0m_tail_outvc1), .B(reset), .Y(s0m_o0sm_n3));
  INV_X0P5B_A12TR s0m_o0sm_u33 (.A(s0m_o0sm_n25), .Y(s0m_o0sm_n35));
  // BSIM@ modules: mx346 
  // BSIM@ covered_modules=1 :   NAND2_X0P5A_A12TR s0m_o0sm_u23 (.A(s0m_o0sm_n24), .B(c0nm_b0m_v0m_n4), .Y(s0m_o0sm_n36));
  NAND3_X0P5A_A12TR s0m_o0sm_u19 (.A(s0m_o0sm_n19), .B(c0nm_b0m_v0m_n4), .C(s0m_o0sm_n21), .Y(s0m_o0sm_n37));
  // BSIM@ modules: mx353 
  // BSIM@ covered_modules=1 :   NOR2_X0P5A_A12TR s0m_o0sm_u14 (.A(reset), .B(s0m_o0sm_n13), .Y(s0m_o0sm_n38));
  AO21A1AI2_X0P5M_A12TR s0m_o0sm_u7 (.A0(s0m_o0sm_n5), .A1(s0m_state_invc1_0_), .B0(s0m_outb1_0_), .C0(s0m_o0sm_n3), .Y(s0m_o0sm_n4));
  NOR2_X0P5A_A12TR s0m_o0sm_u9 (.A(s0m_o0sm_n42), .B(s0m_o0sm_n35), .Y(s0m_o0sm_n41));
  OA21_X0P5M_A12TR s0m_o0sm_u10 (.A0(s0m_o0sm_n6), .A1(s0m_o0sm_n7), .B0(c0nm_b0m_v0m_n4), .Y(s0m_o0sm_n42));
  INV_X0P5B_A12TR s0m_o0sm_u8 (.A(s0m_outb1_1_), .Y(s0m_o0sm_n5));
  // BSIM@ modules: mx272 
  // BSIM@ covered_modules=1 :   NOR3_X0P5A_A12TR s0m_o0sm_u12 (.A(s0m_o0sm_n11), .B(creditin_1), .C(s0m_o0sm_n9), .Y(s0m_o0sm_n6));
  AOI21_X0P5M_A12TR s0m_o0sm_u11 (.A0(creditin_1), .A1(s0m_o0sm_n9), .B0(s0m_n4), .Y(s0m_o0sm_n7));
  NOR3_X0P5A_A12TR s0m_o0sm_u32 (.A(s0m_outb1_1_), .B(s0m_outb1_0_), .C(s0m_debit_outvc1), .Y(s0m_o0sm_n9));
  DFFQ_X1M_A12TR s0m_o0sm_state_assigned_reg (.CK(clk), .Q(s0m_o0sm_state_assigned), .D(s0m_o0sm_n35));
  DFFQ_X1M_A12TR s0m_o0sm_state_credits_reg_0_ (.CK(clk), .Q(s0m_o0sm_state_credits_0_), .D(s0m_o0sm_n36));
  DFFQ_X1M_A12TR s0m_o0sm_state_credits_reg_1_ (.CK(clk), .Q(s0m_o0sm_state_credits_1_), .D(s0m_o0sm_n37));
  DFFQ_X1M_A12TR s0m_o0sm_state_credits_reg_2_ (.CK(clk), .Q(s0m_o0sm_state_credits_2_), .D(s0m_o0sm_n38));
  // BSIM@ modules: mx5 
  // BSIM@ covered_modules=1 :   AOI21_X0P5M_A12TR s0m_m0m_u7 (.A0(s0m_request1[0]), .A1(s0m_m0m_row1_0_), .B0(s0m_m0m_n1), .Y(s0m_outb0_0_));
  OA21_X0P5M_A12TR s0m_m0m_u3 (.A0(s0m_m0m_n1), .A1(s0m_m0m_row1_0_), .B0(s0m_request1[0]), .Y(s0m_outb0_1_));
  AOI21_X0P5M_A12TR s0m_m1m_u7 (.A0(s0m_request1[1]), .A1(s0m_m1m_row1_0_), .B0(s0m_m1m_n1), .Y(s0m_outb1_0_));
  OA21_X0P5M_A12TR s0m_m1m_u3 (.A0(s0m_m1m_n1), .A1(s0m_m1m_row1_0_), .B0(s0m_request1[1]), .Y(s0m_outb1_1_));
  // BSIM@ modules: mx325 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR s0m_u11 (.A(s0m_elig_0_), .B(swalloc_req_0[0]), .Y(s0m_request0[0]));
  // BSIM@ modules: mx324 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR s0m_u10 (.A(s0m_elig_1_), .B(swalloc_req_0[1]), .Y(s0m_request0[1]));
  // BSIM@ modules: mx331 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR s0m_u9 (.A(s0m_elig_0_), .B(swalloc_req_1[0]), .Y(s0m_request1[0]));
  // BSIM@ modules: mx330 
  // BSIM@ covered_modules=1 :   AND2_X0P5M_A12TR s0m_u8 (.A(s0m_elig_1_), .B(swalloc_req_1[1]), .Y(s0m_request1[1]));
  DFFQ_X1M_A12TR s0m_o0nm_state_invc_reg_0_ (.CK(clk), .Q(s0m_state_invc0_0_), .D(s0m_o0nm_n30));
  DFFQ_X1M_A12TR s0m_o0nm_state_invc_reg_1_ (.CK(clk), .Q(s0m_state_invc0_1_), .D(s0m_o0nm_n31));
  DFFQ_X1M_A12TR s0m_o0sm_state_invc_reg_0_ (.CK(clk), .Q(s0m_state_invc1_0_), .D(s0m_o0sm_n27));
  DFFQ_X1M_A12TR s0m_o0sm_state_invc_reg_1_ (.CK(clk), .Q(s0m_state_invc1_1_), .D(s0m_o0sm_n26));
  MXIT2_X0P5M_A12TR s0m_u5 (.A(s0m_n3), .B(s0m_n2), .S0(s0m_state_invc0_0_), .Y(s0m_tail_outvc0));
  // BSIM@ modules: mx26 
  // BSIM@ covered_modules=1 :   MXIT2_X0P5M_A12TR s0m_u3 (.A(s0m_n1), .B(s0m_n2), .S0(s0m_state_invc1_0_), .Y(s0m_tail_outvc1));
  DFFQ_X1M_A12TR c0nm_v0m_state_swreq_reg_0_ (.CK(clk), .Q(swalloc_req_0[0]), .D(c0nm_v0m_n30));
  DFFQ_X1M_A12TR c0nm_v0m_state_swreq_reg_1_ (.CK(clk), .Q(swalloc_req_0[1]), .D(c0nm_v0m_n31));
  DFFQ_X1M_A12TR c0sm_v0m_state_swreq_reg_0_ (.CK(clk), .Q(swalloc_req_1[0]), .D(c0sm_v0m_n33));
  DFFQ_X1M_A12TR c0sm_v0m_state_swreq_reg_1_ (.CK(clk), .Q(swalloc_req_1[1]), .D(c0sm_v0m_n32));
  DFFQ_X1M_A12TR s0m_resp0_reg_0_ (.CK(clk), .Q(swalloc_resp_0[0]), .D(s0m_n25));
  DFFQ_X1M_A12TR s0m_resp0_reg_1_ (.CK(clk), .Q(swalloc_resp_0[1]), .D(s0m_n24));
  DFFQ_X1M_A12TR s0m_resp1_reg_0_ (.CK(clk), .Q(swalloc_resp_1[0]), .D(s0m_n23));
  DFFQ_X1M_A12TR s0m_resp1_reg_1_ (.CK(clk), .Q(swalloc_resp_1[1]), .D(s0m_n22));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_tailout_reg (.CK(clk), .Q(tailout_0), .D(c0nm_b0m_v0m_n1710));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_tailout_reg (.CK(clk), .Q(tailout_1), .D(c0sm_b0m_v0m_n1710));
  TIELO_X1M_A12TR x0m_u3 (.Y(x0m__logic0_));
  // BSIM@ modules: mx341 
  // BSIM@ covered_modules=1 :   TIEHI_X1M_A12TR x0m_u4 (.Y(x0m__logic1_));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx0m_m0m_m0m_u1 (.A(flitout_switch_0[0]), .B(flitout_switch_1[0]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx0m_m0m_int01));
  // BSIM@ modules: mx9 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx0m_m1m_m0m_u1 (.A(flitout_switch_0[0]), .B(flitout_switch_1[0]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx0m_m1m_int01));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx10m_m0m_m0m_u1 (.A(flitout_switch_0[10]), .B(flitout_switch_1[10]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx10m_m0m_int01));
  // BSIM@ modules: mx101 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx10m_m1m_m0m_u1 (.A(flitout_switch_0[10]), .B(flitout_switch_1[10]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx10m_m1m_int01));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx11m_m0m_m0m_u1 (.A(flitout_switch_0[11]), .B(flitout_switch_1[11]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx11m_m0m_int01));
  // BSIM@ modules: mx9 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx11m_m1m_m0m_u1 (.A(flitout_switch_0[11]), .B(flitout_switch_1[11]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx11m_m1m_int01));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx1m_m0m_m0m_u1 (.A(flitout_switch_0[1]), .B(flitout_switch_1[1]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx1m_m0m_int01));
  // BSIM@ modules: mx9 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx1m_m1m_m0m_u1 (.A(flitout_switch_0[1]), .B(flitout_switch_1[1]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx1m_m1m_int01));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx2m_m0m_m0m_u1 (.A(flitout_switch_0[2]), .B(flitout_switch_1[2]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx2m_m0m_int01));
  // BSIM@ modules: mx101 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx2m_m1m_m0m_u1 (.A(flitout_switch_0[2]), .B(flitout_switch_1[2]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx2m_m1m_int01));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx3m_m0m_m0m_u1 (.A(flitout_switch_0[3]), .B(flitout_switch_1[3]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx3m_m0m_int01));
  // BSIM@ modules: mx101 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx3m_m1m_m0m_u1 (.A(flitout_switch_0[3]), .B(flitout_switch_1[3]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx3m_m1m_int01));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx4m_m0m_m0m_u1 (.A(flitout_switch_0[4]), .B(flitout_switch_1[4]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx4m_m0m_int01));
  // BSIM@ modules: mx9 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx4m_m1m_m0m_u1 (.A(flitout_switch_0[4]), .B(flitout_switch_1[4]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx4m_m1m_int01));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx5m_m0m_m0m_u1 (.A(flitout_switch_0[5]), .B(flitout_switch_1[5]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx5m_m0m_int01));
  // BSIM@ modules: mx101 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx5m_m1m_m0m_u1 (.A(flitout_switch_0[5]), .B(flitout_switch_1[5]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx5m_m1m_int01));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx6m_m0m_m0m_u1 (.A(flitout_switch_0[6]), .B(flitout_switch_1[6]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx6m_m0m_int01));
  // BSIM@ modules: mx101 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx6m_m1m_m0m_u1 (.A(flitout_switch_0[6]), .B(flitout_switch_1[6]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx6m_m1m_int01));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx7m_m0m_m0m_u1 (.A(flitout_switch_0[7]), .B(flitout_switch_1[7]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx7m_m0m_int01));
  // BSIM@ modules: mx101 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx7m_m1m_m0m_u1 (.A(flitout_switch_0[7]), .B(flitout_switch_1[7]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx7m_m1m_int01));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx8m_m0m_m0m_u1 (.A(flitout_switch_0[8]), .B(flitout_switch_1[8]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx8m_m0m_int01));
  // BSIM@ modules: mx101 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx8m_m1m_m0m_u1 (.A(flitout_switch_0[8]), .B(flitout_switch_1[8]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx8m_m1m_int01));
  // BSIM@ modules: mx100 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx9m_m0m_m0m_u1 (.A(flitout_switch_0[9]), .B(flitout_switch_1[9]), .S0(x0m_colsel0reg_0_), .Y(x0m_bx9m_m0m_int01));
  // BSIM@ modules: mx101 
  // BSIM@ covered_modules=1 :   MXT2_X0P5M_A12TR x0m_bx9m_m1m_m0m_u1 (.A(flitout_switch_0[9]), .B(flitout_switch_1[9]), .S0(x0m_colsel1reg_0_), .Y(x0m_bx9m_m1m_int01));
  DFFQ_X1M_A12TR x0m_colsel0reg_reg_0_ (.CK(clk), .Q(x0m_colsel0reg_0_), .D(x0m_n3));
  DFFQ_X1M_A12TR x0m_colsel0reg_reg_1_ (.CK(clk), .Q(x0m_colsel0reg_1_), .D(x0m_n4));
  DFFQ_X1M_A12TR x0m_colsel1reg_reg_0_ (.CK(clk), .Q(x0m_colsel1reg_0_), .D(x0m_n5));
  DFFQ_X1M_A12TR x0m_colsel1reg_reg_1_ (.CK(clk), .Q(x0m_colsel1reg_1_), .D(x0m_n6));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   OR2_X0P5M_A12TR x0m_u8 (.A(colsel0[0]), .B(reset), .Y(x0m_n3));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   OR2_X0P5M_A12TR x0m_u7 (.A(colsel0[1]), .B(reset), .Y(x0m_n4));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   OR2_X0P5M_A12TR x0m_u6 (.A(colsel1[0]), .B(reset), .Y(x0m_n5));
  // BSIM@ modules: mx335 
  // BSIM@ covered_modules=1 :   OR2_X0P5M_A12TR x0m_u5 (.A(colsel1[1]), .B(reset), .Y(x0m_n6));
  /*CASIO@<instance>
     <id>mx5</id>
     <module>mux21_mx0</module>
     <compmap>F1:s0m_u2, F2:s0m_m0m_u7, F3:s0m_m0m_u6, F4:s0m_m0m_u5</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21_mx0 mx5(.s0m_m0m_n1(s0m_m0m_n1), .s0m_m0m_row1_0_(s0m_m0m_row1_0_), .s0m_request1_0_(s0m_request1[0]), .s0m_m0m_n2(s0m_m0m_n2), .s0m_m0m_n3(s0m_m0m_n3));
  /*CASIO@<instance>
     <id>mx9</id>
     <module>mux21_mx1</module>
     <compmap>F1:x0m_bx0m_m1m_m0m_u1, F2:x0m_bx1m_m1m_m0m_u1, F3:x0m_bx4m_m1m_m0m_u1, F4:x0m_bx11m_m1m_m0m_u1</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21_mx1 mx9(.flitout_switch_0_0_(flitout_switch_0[0]), .flitout_switch_0_11_(flitout_switch_0[11]), .flitout_switch_0_1_(flitout_switch_0[1]), .flitout_switch_0_4_(flitout_switch_0[4]), .flitout_switch_1_0_(flitout_switch_1[0]), .flitout_switch_1_11_(flitout_switch_1[11]), .flitout_switch_1_1_(flitout_switch_1[1]), .flitout_switch_1_4_(flitout_switch_1[4]), .x0m_colsel1reg_0_(x0m_colsel1reg_0_), .x0m_bx0m_m1m_int01(x0m_bx0m_m1m_int01), .x0m_bx11m_m1m_int01(x0m_bx11m_m1m_int01), .x0m_bx1m_m1m_int01(x0m_bx1m_m1m_int01), .x0m_bx4m_m1m_int01(x0m_bx4m_m1m_int01));
  /*CASIO@<instance>
     <id>mx10</id>
     <module>mux21_mx2</module>
     <compmap>F1:x0m_bx4m_m1m_m4m_u1, F2:x0m_bx11m_m1m_m4m_u1</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21_mx2 mx10(.x0m__logic0_(x0m__logic0_), .x0m_bx11m_m1m_int01(x0m_bx11m_m1m_int01), .x0m_bx4m_m1m_int01(x0m_bx4m_m1m_int01), .x0m_colsel1reg_1_(x0m_colsel1reg_1_), .flitout_1_11_(flitout_1[11]), .flitout_1_4_(flitout_1[4]));
  /*CASIO@<instance>
     <id>mx15</id>
     <module>mux21i_mx3</module>
     <compmap>F1:c0nm_v0m_u7, F2:c0nm_v0m_u4</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_mx3 mx15(.c0nm_routewire_0_(c0nm_routewire[0]), .c0nm_routewire_1_(c0nm_routewire[1]), .c0nm_v0m_n3(c0nm_v0m_n3), .c0nm_v0m_n4(c0nm_v0m_n4), .c0nm_v0m_n7(c0nm_v0m_n7), .c0nm_v0m_n2(c0nm_v0m_n2), .c0nm_v0m_n6(c0nm_v0m_n6));
  /*CASIO@<instance>
     <id>mx16</id>
     <module>mux21i_mx4</module>
     <compmap>F1:c0nm_v0m_u18, F2:c0nm_v0m_u16</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_mx4 mx16(.c0nm_v0m_n18(c0nm_v0m_n18), .c0nm_v0m_n20(c0nm_v0m_n20), .c0nm_v0m_n21(c0nm_v0m_n21), .c0nm_v0m_state_queuelen_0_(c0nm_v0m_state_queuelen_0_), .c0nm_v0m_state_queuelen_1_(c0nm_v0m_state_queuelen_1_), .c0nm_v0m_n15(c0nm_v0m_n15), .c0nm_v0m_n19(c0nm_v0m_n19));
  /*CASIO@<instance>
     <id>mx21</id>
     <module>mux21i_mx5</module>
     <compmap>F1:c0sm_v0m_u7, F2:c0sm_v0m_u4</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_mx5 mx21(.c0sm_routewire_0_(c0sm_routewire[0]), .c0sm_routewire_1_(c0sm_routewire[1]), .c0sm_v0m_n3(c0sm_v0m_n3), .c0sm_v0m_n4(c0sm_v0m_n4), .c0sm_v0m_n7(c0sm_v0m_n7), .c0sm_v0m_n2(c0sm_v0m_n2), .c0sm_v0m_n6(c0sm_v0m_n6));
  /*CASIO@<instance>
     <id>mx22</id>
     <module>mux21i_mx6</module>
     <compmap>F1:c0sm_v0m_u18, F2:c0sm_v0m_u16</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_mx6 mx22(.c0sm_v0m_n18(c0sm_v0m_n18), .c0sm_v0m_n20(c0sm_v0m_n20), .c0sm_v0m_n21(c0sm_v0m_n21), .c0sm_v0m_state_queuelen_0_(c0sm_v0m_state_queuelen_0_), .c0sm_v0m_state_queuelen_1_(c0sm_v0m_state_queuelen_1_), .c0sm_v0m_n15(c0sm_v0m_n15), .c0sm_v0m_n19(c0sm_v0m_n19));
  /*CASIO@<instance>
     <id>mx23</id>
     <module>mux21i_mx7</module>
     <compmap>F1:s0m_u28, F2:s0m_u25</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_mx7 mx23(.s0m_n13(s0m_n13), .s0m_n14(s0m_n14), .s0m_n15(s0m_n15), .s0m_n17(s0m_n17), .s0m_n18(s0m_n18), .s0m_n22(s0m_n22), .s0m_n23(s0m_n23));
  /*CASIO@<instance>
     <id>mx24</id>
     <module>mux21i_mx8</module>
     <compmap>F1:s0m_u19, F2:s0m_u16</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_mx8 mx24(.s0m_n10(s0m_n10), .s0m_n11(s0m_n11), .s0m_n6(s0m_n6), .s0m_n7(s0m_n7), .s0m_n8(s0m_n8), .s0m_n24(s0m_n24), .s0m_n25(s0m_n25));
  /*CASIO@<instance>
     <id>mx25</id>
     <module>mux21i_mx9</module>
     <compmap>F1:s0m_u36, F2:s0m_u13</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_mx9 mx25(.c0nm_v0m_n9(c0nm_v0m_n9), .s0m_n26(s0m_n26), .s0m_n4(s0m_n4), .s0m_n5(s0m_n5), .s0m_state_invc0_0_(s0m_state_invc0_0_), .nomorebufs_0(nomorebufs_0), .s0m_debit_outvc0(s0m_debit_outvc0));
  /*CASIO@<instance>
     <id>mx26</id>
     <module>mux21i_mx10</module>
     <compmap>F1:s0m_u34, F2:s0m_u3</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_mx10 mx26(.c0nm_v0m_n9(c0nm_v0m_n9), .s0m_n1(s0m_n1), .s0m_n2(s0m_n2), .s0m_n20(s0m_n20), .s0m_state_invc1_0_(s0m_state_invc1_0_), .s0m_debit_outvc1(s0m_debit_outvc1), .s0m_tail_outvc1(s0m_tail_outvc1));
  /*CASIO@<instance>
     <id>mx29</id>
     <module>mux21i_aoi22_mx11</module>
     <compmap>F1:c0nm_r0m_u12, F2:c0sm_r0m_u12</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_aoi22_mx11 mx29(.c0nm_r0m_n13(c0nm_r0m_n13), .c0nm_r0m_n14(c0nm_r0m_n14), .c0sm_r0m_n13(c0sm_r0m_n13), .c0sm_r0m_n14(c0sm_r0m_n14), .curry_0_(curry[0]), .curry_1_(curry[1]), .c0nm_r0m_n12(c0nm_r0m_n12), .c0sm_r0m_n12(c0sm_r0m_n12));
  /*CASIO@<instance>
     <id>mx30</id>
     <module>mux21i_aoi22_mx12</module>
     <compmap>F1:c0nm_b0m_v0m_u96, F2:c0nm_b0m_v0m_u89</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_aoi22_mx12 mx30(.c0nm_b0m_n1(c0nm_b0m_n1), .c0nm_b0m_v0m_n114(c0nm_b0m_v0m_n114), .c0nm_b0m_v0m_n119(c0nm_b0m_v0m_n119), .c0nm_b0m_v0m_n125(c0nm_b0m_v0m_n125), .flitin_0_0_(flitin_0[0]), .flitin_0_1_(flitin_0[1]), .c0nm_b0m_v0m_n118(c0nm_b0m_v0m_n118), .c0nm_b0m_v0m_n127(c0nm_b0m_v0m_n127));
  /*CASIO@<instance>
     <id>mx31</id>
     <module>mux21i_aoi22_mx13</module>
     <compmap>F1:c0nm_b0m_v0m_u181, F2:c0nm_b0m_v0m_u160, F3:c0nm_b0m_v0m_u153, F4:c0nm_b0m_v0m_u146, F5:c0nm_b0m_v0m_u139, F6:c0nm_b0m_v0m_u132, F7:c0nm_b0m_v0m_u125, F8:c0nm_b0m_v0m_u118, F9:c0nm_b0m_v0m_u111, F10:c0nm_b0m_v0m_u104</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_aoi22_mx13 mx31(.c0nm_b0m_n1(c0nm_b0m_n1), .c0nm_b0m_v0m_buffers3_10_(c0nm_b0m_v0m_buffers3_10_), .c0nm_b0m_v0m_buffers3_11_(c0nm_b0m_v0m_buffers3_11_), .c0nm_b0m_v0m_buffers3_2_(c0nm_b0m_v0m_buffers3_2_), .c0nm_b0m_v0m_buffers3_3_(c0nm_b0m_v0m_buffers3_3_), .c0nm_b0m_v0m_buffers3_4_(c0nm_b0m_v0m_buffers3_4_), .c0nm_b0m_v0m_buffers3_5_(c0nm_b0m_v0m_buffers3_5_), .c0nm_b0m_v0m_buffers3_6_(c0nm_b0m_v0m_buffers3_6_), .c0nm_b0m_v0m_buffers3_7_(c0nm_b0m_v0m_buffers3_7_), .c0nm_b0m_v0m_buffers3_8_(c0nm_b0m_v0m_buffers3_8_), .c0nm_b0m_v0m_buffers3_9_(c0nm_b0m_v0m_buffers3_9_), .c0nm_b0m_v0m_n128(c0nm_b0m_v0m_n128), .c0nm_b0m_wdata_10_(c0nm_b0m_wdata_10_), .c0nm_b0m_wdata_11_(c0nm_b0m_wdata_11_), .c0nm_b0m_wdata_2_(c0nm_b0m_wdata_2_), .c0nm_b0m_wdata_3_(c0nm_b0m_wdata_3_), .c0nm_b0m_wdata_4_(c0nm_b0m_wdata_4_), .c0nm_b0m_wdata_5_(c0nm_b0m_wdata_5_), .c0nm_b0m_wdata_6_(c0nm_b0m_wdata_6_), .c0nm_b0m_wdata_7_(c0nm_b0m_wdata_7_), .c0nm_b0m_wdata_8_(c0nm_b0m_wdata_8_), .c0nm_b0m_wdata_9_(c0nm_b0m_wdata_9_), .flitin_0_10_(flitin_0[10]), .flitin_0_11_(flitin_0[11]), .flitin_0_2_(flitin_0[2]), .flitin_0_3_(flitin_0[3]), .flitin_0_4_(flitin_0[4]), .flitin_0_5_(flitin_0[5]), .flitin_0_6_(flitin_0[6]), .flitin_0_7_(flitin_0[7]), .flitin_0_8_(flitin_0[8]), .flitin_0_9_(flitin_0[9]), .c0nm_b0m_v0m_n137(c0nm_b0m_v0m_n137), .c0nm_b0m_v0m_n143(c0nm_b0m_v0m_n143), .c0nm_b0m_v0m_n149(c0nm_b0m_v0m_n149), .c0nm_b0m_v0m_n155(c0nm_b0m_v0m_n155), .c0nm_b0m_v0m_n161(c0nm_b0m_v0m_n161), .c0nm_b0m_v0m_n167(c0nm_b0m_v0m_n167), .c0nm_b0m_v0m_n173(c0nm_b0m_v0m_n173), .c0nm_b0m_v0m_n179(c0nm_b0m_v0m_n179), .c0nm_b0m_v0m_n185(c0nm_b0m_v0m_n185), .c0nm_b0m_v0m_n195(c0nm_b0m_v0m_n195));
  /*CASIO@<instance>
     <id>mx42</id>
     <module>mux21i_aoi22_mx14</module>
     <compmap>F1:c0nm_b0m_v0m_u269, F2:c0nm_b0m_v0m_u264, F3:c0nm_b0m_v0m_u241, F4:c0nm_b0m_v0m_u231, F5:c0nm_b0m_v0m_u226</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_aoi22_mx14 mx42(.c0nm_b0m_v0m_buffers0_0_(c0nm_b0m_v0m_buffers0_0_), .c0nm_b0m_v0m_buffers0_1_(c0nm_b0m_v0m_buffers0_1_), .c0nm_b0m_v0m_buffers0_3_(c0nm_b0m_v0m_buffers0_3_), .c0nm_b0m_v0m_buffers0_5_(c0nm_b0m_v0m_buffers0_5_), .c0nm_b0m_v0m_buffers0_6_(c0nm_b0m_v0m_buffers0_6_), .c0nm_b0m_v0m_n114(c0nm_b0m_v0m_n114), .c0nm_b0m_v0m_n125(c0nm_b0m_v0m_n125), .c0nm_b0m_v0m_n141(c0nm_b0m_v0m_n141), .c0nm_b0m_v0m_n153(c0nm_b0m_v0m_n153), .c0nm_b0m_v0m_n159(c0nm_b0m_v0m_n159), .c0nm_b0m_v0m_n192(c0nm_b0m_v0m_n192), .c0nm_b0m_v0m_n193(c0nm_b0m_v0m_n193), .c0nm_b0m_v0m_n268(c0nm_b0m_v0m_n268), .c0nm_b0m_v0m_n269(c0nm_b0m_v0m_n269), .c0nm_b0m_v0m_n271(c0nm_b0m_v0m_n271), .c0nm_b0m_v0m_n275(c0nm_b0m_v0m_n275), .c0nm_b0m_v0m_n276(c0nm_b0m_v0m_n276));
  /*CASIO@<instance>
     <id>mx53</id>
     <module>mux21i_aoi22_mx15</module>
     <compmap>F1:c0nm_b0m_v0m_u184, F2:c0nm_b0m_v0m_u161, F3:c0nm_b0m_v0m_u154, F4:c0nm_b0m_v0m_u147, F5:c0nm_b0m_v0m_u140, F6:c0nm_b0m_v0m_u133, F7:c0nm_b0m_v0m_u126, F8:c0nm_b0m_v0m_u119, F9:c0nm_b0m_v0m_u112, F10:c0nm_b0m_v0m_u105, F11:c0nm_b0m_v0m_u97, F12:c0nm_b0m_v0m_u90</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_aoi22_mx15 mx53(.c0nm_b0m_v0m_buffers0_0_(c0nm_b0m_v0m_buffers0_0_), .c0nm_b0m_v0m_buffers0_10_(c0nm_b0m_v0m_buffers0_10_), .c0nm_b0m_v0m_buffers0_11_(c0nm_b0m_v0m_buffers0_11_), .c0nm_b0m_v0m_buffers0_1_(c0nm_b0m_v0m_buffers0_1_), .c0nm_b0m_v0m_buffers0_2_(c0nm_b0m_v0m_buffers0_2_), .c0nm_b0m_v0m_buffers0_3_(c0nm_b0m_v0m_buffers0_3_), .c0nm_b0m_v0m_buffers0_4_(c0nm_b0m_v0m_buffers0_4_), .c0nm_b0m_v0m_buffers0_5_(c0nm_b0m_v0m_buffers0_5_), .c0nm_b0m_v0m_buffers0_6_(c0nm_b0m_v0m_buffers0_6_), .c0nm_b0m_v0m_buffers0_7_(c0nm_b0m_v0m_buffers0_7_), .c0nm_b0m_v0m_buffers0_8_(c0nm_b0m_v0m_buffers0_8_), .c0nm_b0m_v0m_buffers0_9_(c0nm_b0m_v0m_buffers0_9_), .c0nm_b0m_v0m_buffers2_0_(c0nm_b0m_v0m_buffers2_0_), .c0nm_b0m_v0m_buffers2_10_(c0nm_b0m_v0m_buffers2_10_), .c0nm_b0m_v0m_buffers2_11_(c0nm_b0m_v0m_buffers2_11_), .c0nm_b0m_v0m_buffers2_1_(c0nm_b0m_v0m_buffers2_1_), .c0nm_b0m_v0m_buffers2_2_(c0nm_b0m_v0m_buffers2_2_), .c0nm_b0m_v0m_buffers2_3_(c0nm_b0m_v0m_buffers2_3_), .c0nm_b0m_v0m_buffers2_4_(c0nm_b0m_v0m_buffers2_4_), .c0nm_b0m_v0m_buffers2_5_(c0nm_b0m_v0m_buffers2_5_), .c0nm_b0m_v0m_buffers2_6_(c0nm_b0m_v0m_buffers2_6_), .c0nm_b0m_v0m_buffers2_7_(c0nm_b0m_v0m_buffers2_7_), .c0nm_b0m_v0m_buffers2_8_(c0nm_b0m_v0m_buffers2_8_), .c0nm_b0m_v0m_buffers2_9_(c0nm_b0m_v0m_buffers2_9_), .c0nm_b0m_v0m_n120(c0nm_b0m_v0m_n120), .c0nm_b0m_v0m_n121(c0nm_b0m_v0m_n121), .c0nm_b0m_v0m_n117(c0nm_b0m_v0m_n117), .c0nm_b0m_v0m_n126(c0nm_b0m_v0m_n126), .c0nm_b0m_v0m_n136(c0nm_b0m_v0m_n136), .c0nm_b0m_v0m_n142(c0nm_b0m_v0m_n142), .c0nm_b0m_v0m_n148(c0nm_b0m_v0m_n148), .c0nm_b0m_v0m_n154(c0nm_b0m_v0m_n154), .c0nm_b0m_v0m_n160(c0nm_b0m_v0m_n160), .c0nm_b0m_v0m_n166(c0nm_b0m_v0m_n166), .c0nm_b0m_v0m_n172(c0nm_b0m_v0m_n172), .c0nm_b0m_v0m_n178(c0nm_b0m_v0m_n178), .c0nm_b0m_v0m_n184(c0nm_b0m_v0m_n184), .c0nm_b0m_v0m_n194(c0nm_b0m_v0m_n194));
  /*CASIO@<instance>
     <id>mx64</id>
     <module>mux21i_aoi22_mx16</module>
     <compmap>F1:c0nm_b0m_v0m_u170, F2:c0nm_b0m_v0m_u158, F3:c0nm_b0m_v0m_u151, F4:c0nm_b0m_v0m_u144, F5:c0nm_b0m_v0m_u137, F6:c0nm_b0m_v0m_u130, F7:c0nm_b0m_v0m_u123, F8:c0nm_b0m_v0m_u116, F9:c0nm_b0m_v0m_u109, F10:c0nm_b0m_v0m_u102</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_aoi22_mx16 mx64(.c0nm_b0m_v0m_buffers0_10_(c0nm_b0m_v0m_buffers0_10_), .c0nm_b0m_v0m_buffers0_11_(c0nm_b0m_v0m_buffers0_11_), .c0nm_b0m_v0m_buffers0_2_(c0nm_b0m_v0m_buffers0_2_), .c0nm_b0m_v0m_buffers0_3_(c0nm_b0m_v0m_buffers0_3_), .c0nm_b0m_v0m_buffers0_4_(c0nm_b0m_v0m_buffers0_4_), .c0nm_b0m_v0m_buffers0_5_(c0nm_b0m_v0m_buffers0_5_), .c0nm_b0m_v0m_buffers0_6_(c0nm_b0m_v0m_buffers0_6_), .c0nm_b0m_v0m_buffers0_7_(c0nm_b0m_v0m_buffers0_7_), .c0nm_b0m_v0m_buffers0_8_(c0nm_b0m_v0m_buffers0_8_), .c0nm_b0m_v0m_buffers0_9_(c0nm_b0m_v0m_buffers0_9_), .c0nm_b0m_v0m_n113(c0nm_b0m_v0m_n113), .c0nm_b0m_v0m_n115(c0nm_b0m_v0m_n115), .c0nm_b0m_v0m_n134(c0nm_b0m_v0m_n134), .c0nm_b0m_v0m_n141(c0nm_b0m_v0m_n141), .c0nm_b0m_v0m_n147(c0nm_b0m_v0m_n147), .c0nm_b0m_v0m_n153(c0nm_b0m_v0m_n153), .c0nm_b0m_v0m_n159(c0nm_b0m_v0m_n159), .c0nm_b0m_v0m_n165(c0nm_b0m_v0m_n165), .c0nm_b0m_v0m_n171(c0nm_b0m_v0m_n171), .c0nm_b0m_v0m_n177(c0nm_b0m_v0m_n177), .c0nm_b0m_v0m_n183(c0nm_b0m_v0m_n183), .c0nm_b0m_v0m_n190(c0nm_b0m_v0m_n190), .c0nm_b0m_v0m_n133(c0nm_b0m_v0m_n133), .c0nm_b0m_v0m_n140(c0nm_b0m_v0m_n140), .c0nm_b0m_v0m_n146(c0nm_b0m_v0m_n146), .c0nm_b0m_v0m_n152(c0nm_b0m_v0m_n152), .c0nm_b0m_v0m_n158(c0nm_b0m_v0m_n158), .c0nm_b0m_v0m_n164(c0nm_b0m_v0m_n164), .c0nm_b0m_v0m_n170(c0nm_b0m_v0m_n170), .c0nm_b0m_v0m_n176(c0nm_b0m_v0m_n176), .c0nm_b0m_v0m_n182(c0nm_b0m_v0m_n182), .c0nm_b0m_v0m_n189(c0nm_b0m_v0m_n189));
  /*CASIO@<instance>
     <id>mx65</id>
     <module>mux21i_aoi22_mx17</module>
     <compmap>F1:c0sm_b0m_v0m_u96, F2:c0sm_b0m_v0m_u89</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_aoi22_mx17 mx65(.c0sm_b0m_n2(c0sm_b0m_n2), .c0sm_b0m_v0m_n114(c0sm_b0m_v0m_n114), .c0sm_b0m_v0m_n119(c0sm_b0m_v0m_n119), .c0sm_b0m_v0m_n125(c0sm_b0m_v0m_n125), .flitin_1_0_(flitin_1[0]), .flitin_1_1_(flitin_1[1]), .c0sm_b0m_v0m_n118(c0sm_b0m_v0m_n118), .c0sm_b0m_v0m_n127(c0sm_b0m_v0m_n127));
  /*CASIO@<instance>
     <id>mx66</id>
     <module>mux21i_aoi22_mx18</module>
     <compmap>F1:c0sm_b0m_v0m_u181, F2:c0sm_b0m_v0m_u160, F3:c0sm_b0m_v0m_u153, F4:c0sm_b0m_v0m_u146, F5:c0sm_b0m_v0m_u139, F6:c0sm_b0m_v0m_u132, F7:c0sm_b0m_v0m_u125, F8:c0sm_b0m_v0m_u118, F9:c0sm_b0m_v0m_u111, F10:c0sm_b0m_v0m_u104</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_aoi22_mx18 mx66(.c0sm_b0m_n2(c0sm_b0m_n2), .c0sm_b0m_v0m_buffers3_10_(c0sm_b0m_v0m_buffers3_10_), .c0sm_b0m_v0m_buffers3_11_(c0sm_b0m_v0m_buffers3_11_), .c0sm_b0m_v0m_buffers3_2_(c0sm_b0m_v0m_buffers3_2_), .c0sm_b0m_v0m_buffers3_3_(c0sm_b0m_v0m_buffers3_3_), .c0sm_b0m_v0m_buffers3_4_(c0sm_b0m_v0m_buffers3_4_), .c0sm_b0m_v0m_buffers3_5_(c0sm_b0m_v0m_buffers3_5_), .c0sm_b0m_v0m_buffers3_6_(c0sm_b0m_v0m_buffers3_6_), .c0sm_b0m_v0m_buffers3_7_(c0sm_b0m_v0m_buffers3_7_), .c0sm_b0m_v0m_buffers3_8_(c0sm_b0m_v0m_buffers3_8_), .c0sm_b0m_v0m_buffers3_9_(c0sm_b0m_v0m_buffers3_9_), .c0sm_b0m_v0m_n128(c0sm_b0m_v0m_n128), .c0sm_b0m_wdata_10_(c0sm_b0m_wdata_10_), .c0sm_b0m_wdata_11_(c0sm_b0m_wdata_11_), .c0sm_b0m_wdata_2_(c0sm_b0m_wdata_2_), .c0sm_b0m_wdata_3_(c0sm_b0m_wdata_3_), .c0sm_b0m_wdata_4_(c0sm_b0m_wdata_4_), .c0sm_b0m_wdata_5_(c0sm_b0m_wdata_5_), .c0sm_b0m_wdata_6_(c0sm_b0m_wdata_6_), .c0sm_b0m_wdata_7_(c0sm_b0m_wdata_7_), .c0sm_b0m_wdata_8_(c0sm_b0m_wdata_8_), .c0sm_b0m_wdata_9_(c0sm_b0m_wdata_9_), .flitin_1_10_(flitin_1[10]), .flitin_1_11_(flitin_1[11]), .flitin_1_2_(flitin_1[2]), .flitin_1_3_(flitin_1[3]), .flitin_1_4_(flitin_1[4]), .flitin_1_5_(flitin_1[5]), .flitin_1_6_(flitin_1[6]), .flitin_1_7_(flitin_1[7]), .flitin_1_8_(flitin_1[8]), .flitin_1_9_(flitin_1[9]), .c0sm_b0m_v0m_n137(c0sm_b0m_v0m_n137), .c0sm_b0m_v0m_n143(c0sm_b0m_v0m_n143), .c0sm_b0m_v0m_n149(c0sm_b0m_v0m_n149), .c0sm_b0m_v0m_n155(c0sm_b0m_v0m_n155), .c0sm_b0m_v0m_n161(c0sm_b0m_v0m_n161), .c0sm_b0m_v0m_n167(c0sm_b0m_v0m_n167), .c0sm_b0m_v0m_n173(c0sm_b0m_v0m_n173), .c0sm_b0m_v0m_n179(c0sm_b0m_v0m_n179), .c0sm_b0m_v0m_n185(c0sm_b0m_v0m_n185), .c0sm_b0m_v0m_n195(c0sm_b0m_v0m_n195));
  /*CASIO@<instance>
     <id>mx77</id>
     <module>mux21i_aoi22_mx19</module>
     <compmap>F1:c0sm_b0m_v0m_u241, F2:c0sm_b0m_v0m_u231, F3:c0sm_b0m_v0m_u226</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_aoi22_mx19 mx77(.c0sm_b0m_v0m_buffers0_3_(c0sm_b0m_v0m_buffers0_3_), .c0sm_b0m_v0m_buffers0_5_(c0sm_b0m_v0m_buffers0_5_), .c0sm_b0m_v0m_buffers0_6_(c0sm_b0m_v0m_buffers0_6_), .c0sm_b0m_v0m_n141(c0sm_b0m_v0m_n141), .c0sm_b0m_v0m_n153(c0sm_b0m_v0m_n153), .c0sm_b0m_v0m_n159(c0sm_b0m_v0m_n159), .c0sm_b0m_v0m_n192(c0sm_b0m_v0m_n192), .c0sm_b0m_v0m_n193(c0sm_b0m_v0m_n193), .c0sm_b0m_v0m_n268(c0sm_b0m_v0m_n268), .c0sm_b0m_v0m_n269(c0sm_b0m_v0m_n269), .c0sm_b0m_v0m_n271(c0sm_b0m_v0m_n271));
  /*CASIO@<instance>
     <id>mx88</id>
     <module>mux21i_aoi22_mx20</module>
     <compmap>F1:c0sm_b0m_v0m_u184, F2:c0sm_b0m_v0m_u161, F3:c0sm_b0m_v0m_u154, F4:c0sm_b0m_v0m_u147, F5:c0sm_b0m_v0m_u140, F6:c0sm_b0m_v0m_u133, F7:c0sm_b0m_v0m_u126, F8:c0sm_b0m_v0m_u119, F9:c0sm_b0m_v0m_u112, F10:c0sm_b0m_v0m_u105, F11:c0sm_b0m_v0m_u97, F12:c0sm_b0m_v0m_u90</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_aoi22_mx20 mx88(.c0sm_b0m_v0m_buffers0_0_(c0sm_b0m_v0m_buffers0_0_), .c0sm_b0m_v0m_buffers0_10_(c0sm_b0m_v0m_buffers0_10_), .c0sm_b0m_v0m_buffers0_11_(c0sm_b0m_v0m_buffers0_11_), .c0sm_b0m_v0m_buffers0_1_(c0sm_b0m_v0m_buffers0_1_), .c0sm_b0m_v0m_buffers0_2_(c0sm_b0m_v0m_buffers0_2_), .c0sm_b0m_v0m_buffers0_3_(c0sm_b0m_v0m_buffers0_3_), .c0sm_b0m_v0m_buffers0_4_(c0sm_b0m_v0m_buffers0_4_), .c0sm_b0m_v0m_buffers0_5_(c0sm_b0m_v0m_buffers0_5_), .c0sm_b0m_v0m_buffers0_6_(c0sm_b0m_v0m_buffers0_6_), .c0sm_b0m_v0m_buffers0_7_(c0sm_b0m_v0m_buffers0_7_), .c0sm_b0m_v0m_buffers0_8_(c0sm_b0m_v0m_buffers0_8_), .c0sm_b0m_v0m_buffers0_9_(c0sm_b0m_v0m_buffers0_9_), .c0sm_b0m_v0m_buffers2_0_(c0sm_b0m_v0m_buffers2_0_), .c0sm_b0m_v0m_buffers2_10_(c0sm_b0m_v0m_buffers2_10_), .c0sm_b0m_v0m_buffers2_11_(c0sm_b0m_v0m_buffers2_11_), .c0sm_b0m_v0m_buffers2_1_(c0sm_b0m_v0m_buffers2_1_), .c0sm_b0m_v0m_buffers2_2_(c0sm_b0m_v0m_buffers2_2_), .c0sm_b0m_v0m_buffers2_3_(c0sm_b0m_v0m_buffers2_3_), .c0sm_b0m_v0m_buffers2_4_(c0sm_b0m_v0m_buffers2_4_), .c0sm_b0m_v0m_buffers2_5_(c0sm_b0m_v0m_buffers2_5_), .c0sm_b0m_v0m_buffers2_6_(c0sm_b0m_v0m_buffers2_6_), .c0sm_b0m_v0m_buffers2_7_(c0sm_b0m_v0m_buffers2_7_), .c0sm_b0m_v0m_buffers2_8_(c0sm_b0m_v0m_buffers2_8_), .c0sm_b0m_v0m_buffers2_9_(c0sm_b0m_v0m_buffers2_9_), .c0sm_b0m_v0m_n120(c0sm_b0m_v0m_n120), .c0sm_b0m_v0m_n121(c0sm_b0m_v0m_n121), .c0sm_b0m_v0m_n117(c0sm_b0m_v0m_n117), .c0sm_b0m_v0m_n126(c0sm_b0m_v0m_n126), .c0sm_b0m_v0m_n136(c0sm_b0m_v0m_n136), .c0sm_b0m_v0m_n142(c0sm_b0m_v0m_n142), .c0sm_b0m_v0m_n148(c0sm_b0m_v0m_n148), .c0sm_b0m_v0m_n154(c0sm_b0m_v0m_n154), .c0sm_b0m_v0m_n160(c0sm_b0m_v0m_n160), .c0sm_b0m_v0m_n166(c0sm_b0m_v0m_n166), .c0sm_b0m_v0m_n172(c0sm_b0m_v0m_n172), .c0sm_b0m_v0m_n178(c0sm_b0m_v0m_n178), .c0sm_b0m_v0m_n184(c0sm_b0m_v0m_n184), .c0sm_b0m_v0m_n194(c0sm_b0m_v0m_n194));
  /*CASIO@<instance>
     <id>mx99</id>
     <module>mux21i_aoi22_mx21</module>
     <compmap>F1:c0sm_b0m_v0m_u170, F2:c0sm_b0m_v0m_u158, F3:c0sm_b0m_v0m_u151, F4:c0sm_b0m_v0m_u144, F5:c0sm_b0m_v0m_u137, F6:c0sm_b0m_v0m_u130, F7:c0sm_b0m_v0m_u123, F8:c0sm_b0m_v0m_u116, F9:c0sm_b0m_v0m_u109, F10:c0sm_b0m_v0m_u102</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_aoi22_mx21 mx99(.c0sm_b0m_v0m_buffers0_10_(c0sm_b0m_v0m_buffers0_10_), .c0sm_b0m_v0m_buffers0_11_(c0sm_b0m_v0m_buffers0_11_), .c0sm_b0m_v0m_buffers0_2_(c0sm_b0m_v0m_buffers0_2_), .c0sm_b0m_v0m_buffers0_3_(c0sm_b0m_v0m_buffers0_3_), .c0sm_b0m_v0m_buffers0_4_(c0sm_b0m_v0m_buffers0_4_), .c0sm_b0m_v0m_buffers0_5_(c0sm_b0m_v0m_buffers0_5_), .c0sm_b0m_v0m_buffers0_6_(c0sm_b0m_v0m_buffers0_6_), .c0sm_b0m_v0m_buffers0_7_(c0sm_b0m_v0m_buffers0_7_), .c0sm_b0m_v0m_buffers0_8_(c0sm_b0m_v0m_buffers0_8_), .c0sm_b0m_v0m_buffers0_9_(c0sm_b0m_v0m_buffers0_9_), .c0sm_b0m_v0m_n113(c0sm_b0m_v0m_n113), .c0sm_b0m_v0m_n115(c0sm_b0m_v0m_n115), .c0sm_b0m_v0m_n134(c0sm_b0m_v0m_n134), .c0sm_b0m_v0m_n141(c0sm_b0m_v0m_n141), .c0sm_b0m_v0m_n147(c0sm_b0m_v0m_n147), .c0sm_b0m_v0m_n153(c0sm_b0m_v0m_n153), .c0sm_b0m_v0m_n159(c0sm_b0m_v0m_n159), .c0sm_b0m_v0m_n165(c0sm_b0m_v0m_n165), .c0sm_b0m_v0m_n171(c0sm_b0m_v0m_n171), .c0sm_b0m_v0m_n177(c0sm_b0m_v0m_n177), .c0sm_b0m_v0m_n183(c0sm_b0m_v0m_n183), .c0sm_b0m_v0m_n190(c0sm_b0m_v0m_n190), .c0sm_b0m_v0m_n133(c0sm_b0m_v0m_n133), .c0sm_b0m_v0m_n140(c0sm_b0m_v0m_n140), .c0sm_b0m_v0m_n146(c0sm_b0m_v0m_n146), .c0sm_b0m_v0m_n152(c0sm_b0m_v0m_n152), .c0sm_b0m_v0m_n158(c0sm_b0m_v0m_n158), .c0sm_b0m_v0m_n164(c0sm_b0m_v0m_n164), .c0sm_b0m_v0m_n170(c0sm_b0m_v0m_n170), .c0sm_b0m_v0m_n176(c0sm_b0m_v0m_n176), .c0sm_b0m_v0m_n182(c0sm_b0m_v0m_n182), .c0sm_b0m_v0m_n189(c0sm_b0m_v0m_n189));
  /*CASIO@<instance>
     <id>mx100</id>
     <module>mux31b_mx22</module>
     <compmap>F1:x0m_bx0m_m0m_m0m_u1, F2:x0m_bx0m_m0m_m4m_u1, F3:x0m_bx1m_m0m_m0m_u1, F4:x0m_bx1m_m0m_m4m_u1, F5:x0m_bx2m_m0m_m0m_u1, F6:x0m_bx2m_m0m_m4m_u1, F7:x0m_bx3m_m0m_m0m_u1, F8:x0m_bx3m_m0m_m4m_u1, F9:x0m_bx4m_m0m_m0m_u1, F10:x0m_bx4m_m0m_m4m_u1, F11:x0m_bx5m_m0m_m0m_u1, F12:x0m_bx5m_m0m_m4m_u1, F13:x0m_bx6m_m0m_m0m_u1, F14:x0m_bx6m_m0m_m4m_u1, F15:x0m_bx7m_m0m_m0m_u1, F16:x0m_bx7m_m0m_m4m_u1, F17:x0m_bx8m_m0m_m0m_u1, F18:x0m_bx8m_m0m_m4m_u1, F19:x0m_bx9m_m0m_m0m_u1, F20:x0m_bx9m_m0m_m4m_u1, F21:x0m_bx10m_m0m_m0m_u1, F22:x0m_bx10m_m0m_m4m_u1, F23:x0m_bx11m_m0m_m0m_u1, F24:x0m_bx11m_m0m_m4m_u1</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux31b_mx22 mx100(.flitout_switch_0_0_(flitout_switch_0[0]), .flitout_switch_0_10_(flitout_switch_0[10]), .flitout_switch_0_11_(flitout_switch_0[11]), .flitout_switch_0_1_(flitout_switch_0[1]), .flitout_switch_0_2_(flitout_switch_0[2]), .flitout_switch_0_3_(flitout_switch_0[3]), .flitout_switch_0_4_(flitout_switch_0[4]), .flitout_switch_0_5_(flitout_switch_0[5]), .flitout_switch_0_6_(flitout_switch_0[6]), .flitout_switch_0_7_(flitout_switch_0[7]), .flitout_switch_0_8_(flitout_switch_0[8]), .flitout_switch_0_9_(flitout_switch_0[9]), .flitout_switch_1_0_(flitout_switch_1[0]), .flitout_switch_1_10_(flitout_switch_1[10]), .flitout_switch_1_11_(flitout_switch_1[11]), .flitout_switch_1_1_(flitout_switch_1[1]), .flitout_switch_1_2_(flitout_switch_1[2]), .flitout_switch_1_3_(flitout_switch_1[3]), .flitout_switch_1_4_(flitout_switch_1[4]), .flitout_switch_1_5_(flitout_switch_1[5]), .flitout_switch_1_6_(flitout_switch_1[6]), .flitout_switch_1_7_(flitout_switch_1[7]), .flitout_switch_1_8_(flitout_switch_1[8]), .flitout_switch_1_9_(flitout_switch_1[9]), .x0m__logic0_(x0m__logic0_), .x0m__logic1_(x0m__logic1_), .x0m_colsel0reg_0_(x0m_colsel0reg_0_), .x0m_colsel0reg_1_(x0m_colsel0reg_1_), .flitout_0_0_(flitout_0[0]), .flitout_0_10_(flitout_0[10]), .flitout_0_11_(flitout_0[11]), .flitout_0_1_(flitout_0[1]), .flitout_0_2_(flitout_0[2]), .flitout_0_3_(flitout_0[3]), .flitout_0_4_(flitout_0[4]), .flitout_0_5_(flitout_0[5]), .flitout_0_6_(flitout_0[6]), .flitout_0_7_(flitout_0[7]), .flitout_0_8_(flitout_0[8]), .flitout_0_9_(flitout_0[9]));
  /*CASIO@<instance>
     <id>mx101</id>
     <module>mux31b_mx23</module>
     <compmap>F1:x0m_bx2m_m1m_m0m_u1, F2:x0m_bx2m_m1m_m4m_u1, F3:x0m_bx3m_m1m_m0m_u1, F4:x0m_bx3m_m1m_m4m_u1, F5:x0m_bx5m_m1m_m0m_u1, F6:x0m_bx5m_m1m_m4m_u1, F7:x0m_bx6m_m1m_m0m_u1, F8:x0m_bx6m_m1m_m4m_u1, F9:x0m_bx7m_m1m_m0m_u1, F10:x0m_bx7m_m1m_m4m_u1, F11:x0m_bx8m_m1m_m0m_u1, F12:x0m_bx8m_m1m_m4m_u1, F13:x0m_bx9m_m1m_m0m_u1, F14:x0m_bx9m_m1m_m4m_u1, F15:x0m_bx10m_m1m_m0m_u1, F16:x0m_bx10m_m1m_m4m_u1</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux31b_mx23 mx101(.flitout_switch_0_10_(flitout_switch_0[10]), .flitout_switch_0_2_(flitout_switch_0[2]), .flitout_switch_0_3_(flitout_switch_0[3]), .flitout_switch_0_5_(flitout_switch_0[5]), .flitout_switch_0_6_(flitout_switch_0[6]), .flitout_switch_0_7_(flitout_switch_0[7]), .flitout_switch_0_8_(flitout_switch_0[8]), .flitout_switch_0_9_(flitout_switch_0[9]), .flitout_switch_1_10_(flitout_switch_1[10]), .flitout_switch_1_2_(flitout_switch_1[2]), .flitout_switch_1_3_(flitout_switch_1[3]), .flitout_switch_1_5_(flitout_switch_1[5]), .flitout_switch_1_6_(flitout_switch_1[6]), .flitout_switch_1_7_(flitout_switch_1[7]), .flitout_switch_1_8_(flitout_switch_1[8]), .flitout_switch_1_9_(flitout_switch_1[9]), .x0m__logic0_(x0m__logic0_), .x0m_colsel1reg_0_(x0m_colsel1reg_0_), .x0m_colsel1reg_1_(x0m_colsel1reg_1_), .flitout_1_10_(flitout_1[10]), .flitout_1_2_(flitout_1[2]), .flitout_1_3_(flitout_1[3]), .flitout_1_5_(flitout_1[5]), .flitout_1_6_(flitout_1[6]), .flitout_1_7_(flitout_1[7]), .flitout_1_8_(flitout_1[8]), .flitout_1_9_(flitout_1[9]));
  /*CASIO@<instance>
     <id>mx102</id>
     <module>mux31i_oai222_mx24</module>
     <compmap>F1:c0nm_b0m_v0m_u162, F2:c0nm_b0m_v0m_u155, F3:c0nm_b0m_v0m_u148, F4:c0nm_b0m_v0m_u141, F5:c0nm_b0m_v0m_u134, F6:c0nm_b0m_v0m_u127, F7:c0nm_b0m_v0m_u120, F8:c0nm_b0m_v0m_u113, F9:c0nm_b0m_v0m_u106, F10:c0nm_b0m_v0m_u99</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux31i_oai222_mx24 mx102(.c0nm_b0m_v0m_n107(c0nm_b0m_v0m_n107), .c0nm_b0m_v0m_n129(c0nm_b0m_v0m_n129), .c0nm_b0m_v0m_n130(c0nm_b0m_v0m_n130), .c0nm_b0m_v0m_n131(c0nm_b0m_v0m_n131), .c0nm_b0m_v0m_n138(c0nm_b0m_v0m_n138), .c0nm_b0m_v0m_n144(c0nm_b0m_v0m_n144), .c0nm_b0m_v0m_n150(c0nm_b0m_v0m_n150), .c0nm_b0m_v0m_n156(c0nm_b0m_v0m_n156), .c0nm_b0m_v0m_n162(c0nm_b0m_v0m_n162), .c0nm_b0m_v0m_n168(c0nm_b0m_v0m_n168), .c0nm_b0m_v0m_n17(c0nm_b0m_v0m_n17), .c0nm_b0m_v0m_n174(c0nm_b0m_v0m_n174), .c0nm_b0m_v0m_n180(c0nm_b0m_v0m_n180), .c0nm_b0m_v0m_n186(c0nm_b0m_v0m_n186), .c0nm_b0m_v0m_n19(c0nm_b0m_v0m_n19), .c0nm_b0m_v0m_n33(c0nm_b0m_v0m_n33), .c0nm_b0m_v0m_n34(c0nm_b0m_v0m_n34), .c0nm_b0m_v0m_n36(c0nm_b0m_v0m_n36), .c0nm_b0m_v0m_n37(c0nm_b0m_v0m_n37), .c0nm_b0m_v0m_n39(c0nm_b0m_v0m_n39), .c0nm_b0m_v0m_n40(c0nm_b0m_v0m_n40), .c0nm_b0m_v0m_n42(c0nm_b0m_v0m_n42), .c0nm_b0m_v0m_n43(c0nm_b0m_v0m_n43), .c0nm_b0m_v0m_n45(c0nm_b0m_v0m_n45), .c0nm_b0m_v0m_n46(c0nm_b0m_v0m_n46), .c0nm_b0m_v0m_n48(c0nm_b0m_v0m_n48), .c0nm_b0m_v0m_n49(c0nm_b0m_v0m_n49), .c0nm_b0m_v0m_n63(c0nm_b0m_v0m_n63), .c0nm_b0m_v0m_n64(c0nm_b0m_v0m_n64), .c0nm_b0m_v0m_n66(c0nm_b0m_v0m_n66), .c0nm_b0m_v0m_n67(c0nm_b0m_v0m_n67), .c0nm_b0m_v0m_n69(c0nm_b0m_v0m_n69), .c0nm_b0m_v0m_n70(c0nm_b0m_v0m_n70), .c0nm_b0m_v0m_n208(c0nm_b0m_v0m_n208), .c0nm_b0m_v0m_n209(c0nm_b0m_v0m_n209), .c0nm_b0m_v0m_n210(c0nm_b0m_v0m_n210), .c0nm_b0m_v0m_n211(c0nm_b0m_v0m_n211), .c0nm_b0m_v0m_n212(c0nm_b0m_v0m_n212), .c0nm_b0m_v0m_n213(c0nm_b0m_v0m_n213), .c0nm_b0m_v0m_n214(c0nm_b0m_v0m_n214), .c0nm_b0m_v0m_n215(c0nm_b0m_v0m_n215), .c0nm_b0m_v0m_n216(c0nm_b0m_v0m_n216), .c0nm_b0m_v0m_n217(c0nm_b0m_v0m_n217));
  /*CASIO@<instance>
     <id>mx104</id>
     <module>mux31i_oai222_mx25</module>
     <compmap>F1:c0nm_b0m_v0m_u58, F2:c0nm_b0m_v0m_u56, F3:c0nm_b0m_v0m_u54, F4:c0nm_b0m_v0m_u52, F5:c0nm_b0m_v0m_u50, F6:c0nm_b0m_v0m_u48, F7:c0nm_b0m_v0m_u46, F8:c0nm_b0m_v0m_u44, F9:c0nm_b0m_v0m_u42, F10:c0nm_b0m_v0m_u40</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux31i_oai222_mx25 mx104(.c0nm_b0m_v0m_n17(c0nm_b0m_v0m_n17), .c0nm_b0m_v0m_n19(c0nm_b0m_v0m_n19), .c0nm_b0m_v0m_n33(c0nm_b0m_v0m_n33), .c0nm_b0m_v0m_n34(c0nm_b0m_v0m_n34), .c0nm_b0m_v0m_n36(c0nm_b0m_v0m_n36), .c0nm_b0m_v0m_n37(c0nm_b0m_v0m_n37), .c0nm_b0m_v0m_n39(c0nm_b0m_v0m_n39), .c0nm_b0m_v0m_n40(c0nm_b0m_v0m_n40), .c0nm_b0m_v0m_n42(c0nm_b0m_v0m_n42), .c0nm_b0m_v0m_n43(c0nm_b0m_v0m_n43), .c0nm_b0m_v0m_n45(c0nm_b0m_v0m_n45), .c0nm_b0m_v0m_n46(c0nm_b0m_v0m_n46), .c0nm_b0m_v0m_n48(c0nm_b0m_v0m_n48), .c0nm_b0m_v0m_n49(c0nm_b0m_v0m_n49), .c0nm_b0m_v0m_n63(c0nm_b0m_v0m_n63), .c0nm_b0m_v0m_n64(c0nm_b0m_v0m_n64), .c0nm_b0m_v0m_n66(c0nm_b0m_v0m_n66), .c0nm_b0m_v0m_n67(c0nm_b0m_v0m_n67), .c0nm_b0m_v0m_n69(c0nm_b0m_v0m_n69), .c0nm_b0m_v0m_n70(c0nm_b0m_v0m_n70), .c0nm_b0m_v0m_n76(c0nm_b0m_v0m_n76), .c0nm_b0m_v0m_n81(c0nm_b0m_v0m_n81), .c0nm_b0m_v0m_n82(c0nm_b0m_v0m_n82), .c0nm_b0m_v0m_n83(c0nm_b0m_v0m_n83), .c0nm_b0m_v0m_n84(c0nm_b0m_v0m_n84), .c0nm_b0m_v0m_n85(c0nm_b0m_v0m_n85), .c0nm_b0m_v0m_n86(c0nm_b0m_v0m_n86), .c0nm_b0m_v0m_n87(c0nm_b0m_v0m_n87), .c0nm_b0m_v0m_n88(c0nm_b0m_v0m_n88), .c0nm_b0m_v0m_n89(c0nm_b0m_v0m_n89), .c0nm_b0m_v0m_n90(c0nm_b0m_v0m_n90), .c0nm_b0m_v0m_n91(c0nm_b0m_v0m_n91), .c0nm_b0m_v0m_n92(c0nm_b0m_v0m_n92), .c0nm_b0m_v0m_n232(c0nm_b0m_v0m_n232), .c0nm_b0m_v0m_n233(c0nm_b0m_v0m_n233), .c0nm_b0m_v0m_n234(c0nm_b0m_v0m_n234), .c0nm_b0m_v0m_n235(c0nm_b0m_v0m_n235), .c0nm_b0m_v0m_n236(c0nm_b0m_v0m_n236), .c0nm_b0m_v0m_n237(c0nm_b0m_v0m_n237), .c0nm_b0m_v0m_n238(c0nm_b0m_v0m_n238), .c0nm_b0m_v0m_n239(c0nm_b0m_v0m_n239), .c0nm_b0m_v0m_n240(c0nm_b0m_v0m_n240), .c0nm_b0m_v0m_n241(c0nm_b0m_v0m_n241));
  /*CASIO@<instance>
     <id>mx105</id>
     <module>mux31i_oai222_mx26</module>
     <compmap>F1:c0nm_b0m_v0m_u30, F2:c0nm_b0m_v0m_u29, F3:c0nm_b0m_v0m_u28, F4:c0nm_b0m_v0m_u27, F5:c0nm_b0m_v0m_u26, F6:c0nm_b0m_v0m_u25, F7:c0nm_b0m_v0m_u24, F8:c0nm_b0m_v0m_u23, F9:c0nm_b0m_v0m_u22, F10:c0nm_b0m_v0m_u17</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux31i_oai222_mx26 mx105(.c0nm_b0m_v0m_n17(c0nm_b0m_v0m_n17), .c0nm_b0m_v0m_n18(c0nm_b0m_v0m_n18), .c0nm_b0m_v0m_n19(c0nm_b0m_v0m_n19), .c0nm_b0m_v0m_n20(c0nm_b0m_v0m_n20), .c0nm_b0m_v0m_n21(c0nm_b0m_v0m_n21), .c0nm_b0m_v0m_n22(c0nm_b0m_v0m_n22), .c0nm_b0m_v0m_n33(c0nm_b0m_v0m_n33), .c0nm_b0m_v0m_n34(c0nm_b0m_v0m_n34), .c0nm_b0m_v0m_n35(c0nm_b0m_v0m_n35), .c0nm_b0m_v0m_n36(c0nm_b0m_v0m_n36), .c0nm_b0m_v0m_n37(c0nm_b0m_v0m_n37), .c0nm_b0m_v0m_n38(c0nm_b0m_v0m_n38), .c0nm_b0m_v0m_n39(c0nm_b0m_v0m_n39), .c0nm_b0m_v0m_n40(c0nm_b0m_v0m_n40), .c0nm_b0m_v0m_n41(c0nm_b0m_v0m_n41), .c0nm_b0m_v0m_n42(c0nm_b0m_v0m_n42), .c0nm_b0m_v0m_n43(c0nm_b0m_v0m_n43), .c0nm_b0m_v0m_n44(c0nm_b0m_v0m_n44), .c0nm_b0m_v0m_n45(c0nm_b0m_v0m_n45), .c0nm_b0m_v0m_n46(c0nm_b0m_v0m_n46), .c0nm_b0m_v0m_n47(c0nm_b0m_v0m_n47), .c0nm_b0m_v0m_n48(c0nm_b0m_v0m_n48), .c0nm_b0m_v0m_n49(c0nm_b0m_v0m_n49), .c0nm_b0m_v0m_n62(c0nm_b0m_v0m_n62), .c0nm_b0m_v0m_n63(c0nm_b0m_v0m_n63), .c0nm_b0m_v0m_n64(c0nm_b0m_v0m_n64), .c0nm_b0m_v0m_n65(c0nm_b0m_v0m_n65), .c0nm_b0m_v0m_n66(c0nm_b0m_v0m_n66), .c0nm_b0m_v0m_n67(c0nm_b0m_v0m_n67), .c0nm_b0m_v0m_n68(c0nm_b0m_v0m_n68), .c0nm_b0m_v0m_n69(c0nm_b0m_v0m_n69), .c0nm_b0m_v0m_n70(c0nm_b0m_v0m_n70), .c0nm_b0m_v0m_n71(c0nm_b0m_v0m_n71), .c0nm_b0m_v0m_n244(c0nm_b0m_v0m_n244), .c0nm_b0m_v0m_n245(c0nm_b0m_v0m_n245), .c0nm_b0m_v0m_n246(c0nm_b0m_v0m_n246), .c0nm_b0m_v0m_n247(c0nm_b0m_v0m_n247), .c0nm_b0m_v0m_n248(c0nm_b0m_v0m_n248), .c0nm_b0m_v0m_n249(c0nm_b0m_v0m_n249), .c0nm_b0m_v0m_n250(c0nm_b0m_v0m_n250), .c0nm_b0m_v0m_n251(c0nm_b0m_v0m_n251), .c0nm_b0m_v0m_n252(c0nm_b0m_v0m_n252), .c0nm_b0m_v0m_n255(c0nm_b0m_v0m_n255));
  /*CASIO@<instance>
     <id>mx106</id>
     <module>mux31i_oai222_mx27</module>
     <compmap>F1:c0sm_b0m_v0m_u162, F2:c0sm_b0m_v0m_u155, F3:c0sm_b0m_v0m_u148, F4:c0sm_b0m_v0m_u141, F5:c0sm_b0m_v0m_u134, F6:c0sm_b0m_v0m_u127, F7:c0sm_b0m_v0m_u120, F8:c0sm_b0m_v0m_u113, F9:c0sm_b0m_v0m_u106, F10:c0sm_b0m_v0m_u99</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux31i_oai222_mx27 mx106(.c0sm_b0m_v0m_n107(c0sm_b0m_v0m_n107), .c0sm_b0m_v0m_n129(c0sm_b0m_v0m_n129), .c0sm_b0m_v0m_n130(c0sm_b0m_v0m_n130), .c0sm_b0m_v0m_n131(c0sm_b0m_v0m_n131), .c0sm_b0m_v0m_n138(c0sm_b0m_v0m_n138), .c0sm_b0m_v0m_n144(c0sm_b0m_v0m_n144), .c0sm_b0m_v0m_n150(c0sm_b0m_v0m_n150), .c0sm_b0m_v0m_n156(c0sm_b0m_v0m_n156), .c0sm_b0m_v0m_n162(c0sm_b0m_v0m_n162), .c0sm_b0m_v0m_n168(c0sm_b0m_v0m_n168), .c0sm_b0m_v0m_n17(c0sm_b0m_v0m_n17), .c0sm_b0m_v0m_n174(c0sm_b0m_v0m_n174), .c0sm_b0m_v0m_n180(c0sm_b0m_v0m_n180), .c0sm_b0m_v0m_n186(c0sm_b0m_v0m_n186), .c0sm_b0m_v0m_n19(c0sm_b0m_v0m_n19), .c0sm_b0m_v0m_n33(c0sm_b0m_v0m_n33), .c0sm_b0m_v0m_n34(c0sm_b0m_v0m_n34), .c0sm_b0m_v0m_n36(c0sm_b0m_v0m_n36), .c0sm_b0m_v0m_n37(c0sm_b0m_v0m_n37), .c0sm_b0m_v0m_n39(c0sm_b0m_v0m_n39), .c0sm_b0m_v0m_n40(c0sm_b0m_v0m_n40), .c0sm_b0m_v0m_n42(c0sm_b0m_v0m_n42), .c0sm_b0m_v0m_n43(c0sm_b0m_v0m_n43), .c0sm_b0m_v0m_n45(c0sm_b0m_v0m_n45), .c0sm_b0m_v0m_n46(c0sm_b0m_v0m_n46), .c0sm_b0m_v0m_n48(c0sm_b0m_v0m_n48), .c0sm_b0m_v0m_n49(c0sm_b0m_v0m_n49), .c0sm_b0m_v0m_n63(c0sm_b0m_v0m_n63), .c0sm_b0m_v0m_n64(c0sm_b0m_v0m_n64), .c0sm_b0m_v0m_n66(c0sm_b0m_v0m_n66), .c0sm_b0m_v0m_n67(c0sm_b0m_v0m_n67), .c0sm_b0m_v0m_n69(c0sm_b0m_v0m_n69), .c0sm_b0m_v0m_n70(c0sm_b0m_v0m_n70), .c0sm_b0m_v0m_n321(c0sm_b0m_v0m_n321), .c0sm_b0m_v0m_n322(c0sm_b0m_v0m_n322), .c0sm_b0m_v0m_n323(c0sm_b0m_v0m_n323), .c0sm_b0m_v0m_n324(c0sm_b0m_v0m_n324), .c0sm_b0m_v0m_n325(c0sm_b0m_v0m_n325), .c0sm_b0m_v0m_n326(c0sm_b0m_v0m_n326), .c0sm_b0m_v0m_n327(c0sm_b0m_v0m_n327), .c0sm_b0m_v0m_n328(c0sm_b0m_v0m_n328), .c0sm_b0m_v0m_n329(c0sm_b0m_v0m_n329), .c0sm_b0m_v0m_n330(c0sm_b0m_v0m_n330));
  /*CASIO@<instance>
     <id>mx108</id>
     <module>mux31i_oai222_mx28</module>
     <compmap>F1:c0sm_b0m_v0m_u58, F2:c0sm_b0m_v0m_u56, F3:c0sm_b0m_v0m_u54, F4:c0sm_b0m_v0m_u52, F5:c0sm_b0m_v0m_u50, F6:c0sm_b0m_v0m_u48, F7:c0sm_b0m_v0m_u46, F8:c0sm_b0m_v0m_u44, F9:c0sm_b0m_v0m_u42, F10:c0sm_b0m_v0m_u40</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux31i_oai222_mx28 mx108(.c0sm_b0m_v0m_n17(c0sm_b0m_v0m_n17), .c0sm_b0m_v0m_n19(c0sm_b0m_v0m_n19), .c0sm_b0m_v0m_n33(c0sm_b0m_v0m_n33), .c0sm_b0m_v0m_n34(c0sm_b0m_v0m_n34), .c0sm_b0m_v0m_n36(c0sm_b0m_v0m_n36), .c0sm_b0m_v0m_n37(c0sm_b0m_v0m_n37), .c0sm_b0m_v0m_n39(c0sm_b0m_v0m_n39), .c0sm_b0m_v0m_n40(c0sm_b0m_v0m_n40), .c0sm_b0m_v0m_n42(c0sm_b0m_v0m_n42), .c0sm_b0m_v0m_n43(c0sm_b0m_v0m_n43), .c0sm_b0m_v0m_n45(c0sm_b0m_v0m_n45), .c0sm_b0m_v0m_n46(c0sm_b0m_v0m_n46), .c0sm_b0m_v0m_n48(c0sm_b0m_v0m_n48), .c0sm_b0m_v0m_n49(c0sm_b0m_v0m_n49), .c0sm_b0m_v0m_n63(c0sm_b0m_v0m_n63), .c0sm_b0m_v0m_n64(c0sm_b0m_v0m_n64), .c0sm_b0m_v0m_n66(c0sm_b0m_v0m_n66), .c0sm_b0m_v0m_n67(c0sm_b0m_v0m_n67), .c0sm_b0m_v0m_n69(c0sm_b0m_v0m_n69), .c0sm_b0m_v0m_n70(c0sm_b0m_v0m_n70), .c0sm_b0m_v0m_n76(c0sm_b0m_v0m_n76), .c0sm_b0m_v0m_n81(c0sm_b0m_v0m_n81), .c0sm_b0m_v0m_n82(c0sm_b0m_v0m_n82), .c0sm_b0m_v0m_n83(c0sm_b0m_v0m_n83), .c0sm_b0m_v0m_n84(c0sm_b0m_v0m_n84), .c0sm_b0m_v0m_n85(c0sm_b0m_v0m_n85), .c0sm_b0m_v0m_n86(c0sm_b0m_v0m_n86), .c0sm_b0m_v0m_n87(c0sm_b0m_v0m_n87), .c0sm_b0m_v0m_n88(c0sm_b0m_v0m_n88), .c0sm_b0m_v0m_n89(c0sm_b0m_v0m_n89), .c0sm_b0m_v0m_n90(c0sm_b0m_v0m_n90), .c0sm_b0m_v0m_n91(c0sm_b0m_v0m_n91), .c0sm_b0m_v0m_n92(c0sm_b0m_v0m_n92), .c0sm_b0m_v0m_n297(c0sm_b0m_v0m_n297), .c0sm_b0m_v0m_n298(c0sm_b0m_v0m_n298), .c0sm_b0m_v0m_n299(c0sm_b0m_v0m_n299), .c0sm_b0m_v0m_n300(c0sm_b0m_v0m_n300), .c0sm_b0m_v0m_n301(c0sm_b0m_v0m_n301), .c0sm_b0m_v0m_n302(c0sm_b0m_v0m_n302), .c0sm_b0m_v0m_n303(c0sm_b0m_v0m_n303), .c0sm_b0m_v0m_n304(c0sm_b0m_v0m_n304), .c0sm_b0m_v0m_n305(c0sm_b0m_v0m_n305), .c0sm_b0m_v0m_n306(c0sm_b0m_v0m_n306));
  /*CASIO@<instance>
     <id>mx109</id>
     <module>mux31i_oai222_mx29</module>
     <compmap>F1:c0sm_b0m_v0m_u30, F2:c0sm_b0m_v0m_u29, F3:c0sm_b0m_v0m_u28, F4:c0sm_b0m_v0m_u27, F5:c0sm_b0m_v0m_u26, F6:c0sm_b0m_v0m_u25, F7:c0sm_b0m_v0m_u24, F8:c0sm_b0m_v0m_u23, F9:c0sm_b0m_v0m_u22, F10:c0sm_b0m_v0m_u17</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux31i_oai222_mx29 mx109(.c0sm_b0m_v0m_n17(c0sm_b0m_v0m_n17), .c0sm_b0m_v0m_n18(c0sm_b0m_v0m_n18), .c0sm_b0m_v0m_n19(c0sm_b0m_v0m_n19), .c0sm_b0m_v0m_n20(c0sm_b0m_v0m_n20), .c0sm_b0m_v0m_n21(c0sm_b0m_v0m_n21), .c0sm_b0m_v0m_n22(c0sm_b0m_v0m_n22), .c0sm_b0m_v0m_n33(c0sm_b0m_v0m_n33), .c0sm_b0m_v0m_n34(c0sm_b0m_v0m_n34), .c0sm_b0m_v0m_n35(c0sm_b0m_v0m_n35), .c0sm_b0m_v0m_n36(c0sm_b0m_v0m_n36), .c0sm_b0m_v0m_n37(c0sm_b0m_v0m_n37), .c0sm_b0m_v0m_n38(c0sm_b0m_v0m_n38), .c0sm_b0m_v0m_n39(c0sm_b0m_v0m_n39), .c0sm_b0m_v0m_n40(c0sm_b0m_v0m_n40), .c0sm_b0m_v0m_n41(c0sm_b0m_v0m_n41), .c0sm_b0m_v0m_n42(c0sm_b0m_v0m_n42), .c0sm_b0m_v0m_n43(c0sm_b0m_v0m_n43), .c0sm_b0m_v0m_n44(c0sm_b0m_v0m_n44), .c0sm_b0m_v0m_n45(c0sm_b0m_v0m_n45), .c0sm_b0m_v0m_n46(c0sm_b0m_v0m_n46), .c0sm_b0m_v0m_n47(c0sm_b0m_v0m_n47), .c0sm_b0m_v0m_n48(c0sm_b0m_v0m_n48), .c0sm_b0m_v0m_n49(c0sm_b0m_v0m_n49), .c0sm_b0m_v0m_n62(c0sm_b0m_v0m_n62), .c0sm_b0m_v0m_n63(c0sm_b0m_v0m_n63), .c0sm_b0m_v0m_n64(c0sm_b0m_v0m_n64), .c0sm_b0m_v0m_n65(c0sm_b0m_v0m_n65), .c0sm_b0m_v0m_n66(c0sm_b0m_v0m_n66), .c0sm_b0m_v0m_n67(c0sm_b0m_v0m_n67), .c0sm_b0m_v0m_n68(c0sm_b0m_v0m_n68), .c0sm_b0m_v0m_n69(c0sm_b0m_v0m_n69), .c0sm_b0m_v0m_n70(c0sm_b0m_v0m_n70), .c0sm_b0m_v0m_n71(c0sm_b0m_v0m_n71), .c0sm_b0m_v0m_n283(c0sm_b0m_v0m_n283), .c0sm_b0m_v0m_n286(c0sm_b0m_v0m_n286), .c0sm_b0m_v0m_n287(c0sm_b0m_v0m_n287), .c0sm_b0m_v0m_n288(c0sm_b0m_v0m_n288), .c0sm_b0m_v0m_n289(c0sm_b0m_v0m_n289), .c0sm_b0m_v0m_n290(c0sm_b0m_v0m_n290), .c0sm_b0m_v0m_n291(c0sm_b0m_v0m_n291), .c0sm_b0m_v0m_n292(c0sm_b0m_v0m_n292), .c0sm_b0m_v0m_n293(c0sm_b0m_v0m_n293), .c0sm_b0m_v0m_n294(c0sm_b0m_v0m_n294));
  /*CASIO@<instance>
     <id>mx110</id>
     <module>mux21i_aoi221_mx30</module>
     <compmap>F1:c0nm_r0m_u9, F2:c0sm_r0m_u9</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_aoi221_mx30 mx110(.c0nm_r0m_n10(c0nm_r0m_n10), .c0nm_r0m_n8(c0nm_r0m_n8), .c0nm_r0m_n9(c0nm_r0m_n9), .c0sm_r0m_n10(c0sm_r0m_n10), .c0sm_r0m_n8(c0sm_r0m_n8), .c0sm_r0m_n9(c0sm_r0m_n9), .currx_0_(currx[0]), .currx_1_(currx[1]), .c0nm_r0m_n7(c0nm_r0m_n7), .c0sm_r0m_n7(c0sm_r0m_n7));
  /*CASIO@<instance>
     <id>mx132</id>
     <module>mux21i_aoi221_mx31</module>
     <compmap>F1:c0sm_b0m_v0m_u68, F2:c0sm_b0m_v0m_u66</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_aoi221_mx31 mx132(.c0sm_b0m_v0m_n100(c0sm_b0m_v0m_n100), .c0sm_b0m_v0m_n25(c0sm_b0m_v0m_n25), .c0sm_b0m_v0m_n27(c0sm_b0m_v0m_n27), .c0sm_b0m_v0m_n31(c0sm_b0m_v0m_n31), .c0sm_b0m_v0m_n32(c0sm_b0m_v0m_n32), .c0sm_b0m_v0m_n99(c0sm_b0m_v0m_n99), .reset(reset), .c0sm_b0m_v0m_n101(c0sm_b0m_v0m_n101), .c0sm_b0m_v0m_n97(c0sm_b0m_v0m_n97));
  /*CASIO@<instance>
     <id>mx167</id>
     <module>mux21i_aoi221_mx32</module>
     <compmap>F1:c0nm_b0m_v0m_u68, F2:c0nm_b0m_v0m_u66</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_aoi221_mx32 mx167(.c0nm_b0m_v0m_n100(c0nm_b0m_v0m_n100), .c0nm_b0m_v0m_n25(c0nm_b0m_v0m_n25), .c0nm_b0m_v0m_n27(c0nm_b0m_v0m_n27), .c0nm_b0m_v0m_n31(c0nm_b0m_v0m_n31), .c0nm_b0m_v0m_n32(c0nm_b0m_v0m_n32), .c0nm_b0m_v0m_n99(c0nm_b0m_v0m_n99), .reset(reset), .c0nm_b0m_v0m_n101(c0nm_b0m_v0m_n101), .c0nm_b0m_v0m_n97(c0nm_b0m_v0m_n97));
  /*CASIO@<instance>
     <id>mx194</id>
     <module>mux21i_aoi221_mx33</module>
     <compmap>F1:c0sm_b0m_v0m_u94, F2:c0sm_b0m_v0m_u87</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_aoi221_mx33 mx194(.c0sm_b0m_v0m_buffers0_0_(c0sm_b0m_v0m_buffers0_0_), .c0sm_b0m_v0m_buffers0_1_(c0sm_b0m_v0m_buffers0_1_), .c0sm_b0m_v0m_n113(c0sm_b0m_v0m_n113), .c0sm_b0m_v0m_n114(c0sm_b0m_v0m_n114), .c0sm_b0m_v0m_n115(c0sm_b0m_v0m_n115), .c0sm_b0m_v0m_n125(c0sm_b0m_v0m_n125), .debitout_1(debitout_1), .c0sm_b0m_v0m_n112(c0sm_b0m_v0m_n112), .c0sm_b0m_v0m_n124(c0sm_b0m_v0m_n124));
  /*CASIO@<instance>
     <id>mx207</id>
     <module>mux21_oa221_mx34</module>
     <compmap>F1:c0nm_b0m_v0m_u240, F2:c0nm_b0m_v0m_u230, F3:c0nm_b0m_v0m_u225, F4:c0nm_r0m_u19, F5:c0nm_r0m_u17, F6:c0nm_r0m_u13</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21_oa221_mx34 mx207(.c0nm_b0m_v0m_n138(c0nm_b0m_v0m_n138), .c0nm_b0m_v0m_n150(c0nm_b0m_v0m_n150), .c0nm_b0m_v0m_n156(c0nm_b0m_v0m_n156), .c0nm_b0m_v0m_n187(c0nm_b0m_v0m_n187), .c0nm_b0m_v0m_n268(c0nm_b0m_v0m_n268), .c0nm_b0m_v0m_n269(c0nm_b0m_v0m_n269), .c0nm_b0m_v0m_n271(c0nm_b0m_v0m_n271), .c0nm_b0m_v0m_n38(c0nm_b0m_v0m_n38), .c0nm_b0m_v0m_n44(c0nm_b0m_v0m_n44), .c0nm_b0m_v0m_n47(c0nm_b0m_v0m_n47), .c0nm_b0m_v0m_n73(c0nm_b0m_v0m_n73), .c0nm_r0m_n14(c0nm_r0m_n14), .c0nm_r0m_n8(c0nm_r0m_n8), .c0nm_r0m_n9(c0nm_r0m_n9));
  /*CASIO@<instance>
     <id>mx211</id>
     <module>mux21_oa221_mx35</module>
     <compmap>F1:c0nm_b0m_v0m_u169, F2:c0nm_b0m_v0m_u168, F3:c0nm_b0m_v0m_u157, F4:c0nm_b0m_v0m_u156, F5:c0nm_b0m_v0m_u150, F6:c0nm_b0m_v0m_u149, F7:c0nm_b0m_v0m_u143, F8:c0nm_b0m_v0m_u142, F9:c0nm_b0m_v0m_u136, F10:c0nm_b0m_v0m_u135, F11:c0nm_b0m_v0m_u129, F12:c0nm_b0m_v0m_u128, F13:c0nm_b0m_v0m_u122, F14:c0nm_b0m_v0m_u121, F15:c0nm_b0m_v0m_u115, F16:c0nm_b0m_v0m_u114, F17:c0nm_b0m_v0m_u108, F18:c0nm_b0m_v0m_u107, F19:c0nm_b0m_v0m_u101, F20:c0nm_b0m_v0m_u100</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21_oa221_mx35 mx211(.c0nm_b0m_v0m_n110(c0nm_b0m_v0m_n110), .c0nm_b0m_v0m_n111(c0nm_b0m_v0m_n111), .c0nm_b0m_v0m_n131(c0nm_b0m_v0m_n131), .c0nm_b0m_v0m_n133(c0nm_b0m_v0m_n133), .c0nm_b0m_v0m_n138(c0nm_b0m_v0m_n138), .c0nm_b0m_v0m_n140(c0nm_b0m_v0m_n140), .c0nm_b0m_v0m_n144(c0nm_b0m_v0m_n144), .c0nm_b0m_v0m_n146(c0nm_b0m_v0m_n146), .c0nm_b0m_v0m_n150(c0nm_b0m_v0m_n150), .c0nm_b0m_v0m_n152(c0nm_b0m_v0m_n152), .c0nm_b0m_v0m_n156(c0nm_b0m_v0m_n156), .c0nm_b0m_v0m_n158(c0nm_b0m_v0m_n158), .c0nm_b0m_v0m_n162(c0nm_b0m_v0m_n162), .c0nm_b0m_v0m_n164(c0nm_b0m_v0m_n164), .c0nm_b0m_v0m_n168(c0nm_b0m_v0m_n168), .c0nm_b0m_v0m_n170(c0nm_b0m_v0m_n170), .c0nm_b0m_v0m_n174(c0nm_b0m_v0m_n174), .c0nm_b0m_v0m_n176(c0nm_b0m_v0m_n176), .c0nm_b0m_v0m_n180(c0nm_b0m_v0m_n180), .c0nm_b0m_v0m_n182(c0nm_b0m_v0m_n182), .c0nm_b0m_v0m_n186(c0nm_b0m_v0m_n186), .c0nm_b0m_v0m_n189(c0nm_b0m_v0m_n189), .c0nm_b0m_v0m_n21(c0nm_b0m_v0m_n21), .c0nm_b0m_v0m_n35(c0nm_b0m_v0m_n35), .c0nm_b0m_v0m_n38(c0nm_b0m_v0m_n38), .c0nm_b0m_v0m_n41(c0nm_b0m_v0m_n41), .c0nm_b0m_v0m_n44(c0nm_b0m_v0m_n44), .c0nm_b0m_v0m_n47(c0nm_b0m_v0m_n47), .c0nm_b0m_v0m_n62(c0nm_b0m_v0m_n62), .c0nm_b0m_v0m_n65(c0nm_b0m_v0m_n65), .c0nm_b0m_v0m_n68(c0nm_b0m_v0m_n68), .c0nm_b0m_v0m_n71(c0nm_b0m_v0m_n71), .c0nm_b0m_v0m_n17(c0nm_b0m_v0m_n17), .c0nm_b0m_v0m_n33(c0nm_b0m_v0m_n33), .c0nm_b0m_v0m_n36(c0nm_b0m_v0m_n36), .c0nm_b0m_v0m_n39(c0nm_b0m_v0m_n39), .c0nm_b0m_v0m_n42(c0nm_b0m_v0m_n42), .c0nm_b0m_v0m_n45(c0nm_b0m_v0m_n45), .c0nm_b0m_v0m_n48(c0nm_b0m_v0m_n48), .c0nm_b0m_v0m_n63(c0nm_b0m_v0m_n63), .c0nm_b0m_v0m_n66(c0nm_b0m_v0m_n66), .c0nm_b0m_v0m_n69(c0nm_b0m_v0m_n69));
  /*CASIO@<instance>
     <id>mx212</id>
     <module>mux21_oa221_mx36</module>
     <compmap>F1:c0sm_b0m_v0m_u240, F2:c0sm_b0m_v0m_u230, F3:c0sm_b0m_v0m_u225, F4:c0sm_r0m_u19, F5:c0sm_r0m_u17, F6:c0sm_r0m_u13</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21_oa221_mx36 mx212(.c0sm_b0m_v0m_n138(c0sm_b0m_v0m_n138), .c0sm_b0m_v0m_n150(c0sm_b0m_v0m_n150), .c0sm_b0m_v0m_n156(c0sm_b0m_v0m_n156), .c0sm_b0m_v0m_n187(c0sm_b0m_v0m_n187), .c0sm_b0m_v0m_n268(c0sm_b0m_v0m_n268), .c0sm_b0m_v0m_n269(c0sm_b0m_v0m_n269), .c0sm_b0m_v0m_n271(c0sm_b0m_v0m_n271), .c0sm_b0m_v0m_n38(c0sm_b0m_v0m_n38), .c0sm_b0m_v0m_n44(c0sm_b0m_v0m_n44), .c0sm_b0m_v0m_n47(c0sm_b0m_v0m_n47), .c0sm_b0m_v0m_n73(c0sm_b0m_v0m_n73), .c0sm_r0m_n14(c0sm_r0m_n14), .c0sm_r0m_n8(c0sm_r0m_n8), .c0sm_r0m_n9(c0sm_r0m_n9));
  /*CASIO@<instance>
     <id>mx216</id>
     <module>mux21_oa221_mx37</module>
     <compmap>F1:c0sm_b0m_v0m_u169, F2:c0sm_b0m_v0m_u168, F3:c0sm_b0m_v0m_u157, F4:c0sm_b0m_v0m_u156, F5:c0sm_b0m_v0m_u150, F6:c0sm_b0m_v0m_u149, F7:c0sm_b0m_v0m_u143, F8:c0sm_b0m_v0m_u142, F9:c0sm_b0m_v0m_u136, F10:c0sm_b0m_v0m_u135, F11:c0sm_b0m_v0m_u129, F12:c0sm_b0m_v0m_u128, F13:c0sm_b0m_v0m_u122, F14:c0sm_b0m_v0m_u121, F15:c0sm_b0m_v0m_u115, F16:c0sm_b0m_v0m_u114, F17:c0sm_b0m_v0m_u108, F18:c0sm_b0m_v0m_u107, F19:c0sm_b0m_v0m_u101, F20:c0sm_b0m_v0m_u100</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21_oa221_mx37 mx216(.c0sm_b0m_v0m_n110(c0sm_b0m_v0m_n110), .c0sm_b0m_v0m_n111(c0sm_b0m_v0m_n111), .c0sm_b0m_v0m_n131(c0sm_b0m_v0m_n131), .c0sm_b0m_v0m_n133(c0sm_b0m_v0m_n133), .c0sm_b0m_v0m_n138(c0sm_b0m_v0m_n138), .c0sm_b0m_v0m_n140(c0sm_b0m_v0m_n140), .c0sm_b0m_v0m_n144(c0sm_b0m_v0m_n144), .c0sm_b0m_v0m_n146(c0sm_b0m_v0m_n146), .c0sm_b0m_v0m_n150(c0sm_b0m_v0m_n150), .c0sm_b0m_v0m_n152(c0sm_b0m_v0m_n152), .c0sm_b0m_v0m_n156(c0sm_b0m_v0m_n156), .c0sm_b0m_v0m_n158(c0sm_b0m_v0m_n158), .c0sm_b0m_v0m_n162(c0sm_b0m_v0m_n162), .c0sm_b0m_v0m_n164(c0sm_b0m_v0m_n164), .c0sm_b0m_v0m_n168(c0sm_b0m_v0m_n168), .c0sm_b0m_v0m_n170(c0sm_b0m_v0m_n170), .c0sm_b0m_v0m_n174(c0sm_b0m_v0m_n174), .c0sm_b0m_v0m_n176(c0sm_b0m_v0m_n176), .c0sm_b0m_v0m_n180(c0sm_b0m_v0m_n180), .c0sm_b0m_v0m_n182(c0sm_b0m_v0m_n182), .c0sm_b0m_v0m_n186(c0sm_b0m_v0m_n186), .c0sm_b0m_v0m_n189(c0sm_b0m_v0m_n189), .c0sm_b0m_v0m_n21(c0sm_b0m_v0m_n21), .c0sm_b0m_v0m_n35(c0sm_b0m_v0m_n35), .c0sm_b0m_v0m_n38(c0sm_b0m_v0m_n38), .c0sm_b0m_v0m_n41(c0sm_b0m_v0m_n41), .c0sm_b0m_v0m_n44(c0sm_b0m_v0m_n44), .c0sm_b0m_v0m_n47(c0sm_b0m_v0m_n47), .c0sm_b0m_v0m_n62(c0sm_b0m_v0m_n62), .c0sm_b0m_v0m_n65(c0sm_b0m_v0m_n65), .c0sm_b0m_v0m_n68(c0sm_b0m_v0m_n68), .c0sm_b0m_v0m_n71(c0sm_b0m_v0m_n71), .c0sm_b0m_v0m_n17(c0sm_b0m_v0m_n17), .c0sm_b0m_v0m_n33(c0sm_b0m_v0m_n33), .c0sm_b0m_v0m_n36(c0sm_b0m_v0m_n36), .c0sm_b0m_v0m_n39(c0sm_b0m_v0m_n39), .c0sm_b0m_v0m_n42(c0sm_b0m_v0m_n42), .c0sm_b0m_v0m_n45(c0sm_b0m_v0m_n45), .c0sm_b0m_v0m_n48(c0sm_b0m_v0m_n48), .c0sm_b0m_v0m_n63(c0sm_b0m_v0m_n63), .c0sm_b0m_v0m_n66(c0sm_b0m_v0m_n66), .c0sm_b0m_v0m_n69(c0sm_b0m_v0m_n69));
  /*CASIO@<instance>
     <id>mx244</id>
     <module>mux21i_oai221_mx38</module>
     <compmap>F1:c0sm_b0m_v0m_u93, F2:c0sm_b0m_v0m_u86</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux21i_oai221_mx38 mx244(.c0sm_b0m_v0m_n105(c0sm_b0m_v0m_n105), .c0sm_b0m_v0m_n110(c0sm_b0m_v0m_n110), .c0sm_b0m_v0m_n111(c0sm_b0m_v0m_n111), .c0sm_b0m_v0m_n112(c0sm_b0m_v0m_n112), .c0sm_b0m_v0m_n122(c0sm_b0m_v0m_n122), .c0sm_b0m_v0m_n124(c0sm_b0m_v0m_n124), .c0sm_b0m_v0m_n23(c0sm_b0m_v0m_n23), .c0sm_b0m_v0m_n29(c0sm_b0m_v0m_n29), .c0sm_b0m_v0m_n27(c0sm_b0m_v0m_n27), .c0sm_b0m_v0m_n32(c0sm_b0m_v0m_n32));
  /*CASIO@<instance>
     <id>mx245</id>
     <module>reg_mx39</module>
     <compmap>F1:c0nm_b0m_v0m_u196, F2:c0nm_b0m_v0m_u194, F3:c0nm_b0m_v0m_rdata_reg_0_, F4:c0nm_b0m_v0m_rdata_reg_1_, </compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  reg_mx39 mx245(.c0nm_b0m_v0m_n11(c0nm_b0m_v0m_n11), .c0nm_b0m_v0m_n262(c0nm_b0m_v0m_n262), .c0nm_b0m_v0m_n263(c0nm_b0m_v0m_n263), .clk(clk), .c0nm_b0m_rdata_0_(c0nm_b0m_rdata[0]), .c0nm_b0m_rdata_1_(c0nm_b0m_rdata[1]));
  /*CASIO@<instance>
     <id>mx246</id>
     <module>reg_mx40</module>
     <compmap>F1:c0sm_b0m_v0m_u196, F2:c0sm_b0m_v0m_u194, F3:c0sm_b0m_v0m_rdata_reg_0_, F4:c0sm_b0m_v0m_rdata_reg_1_, </compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  reg_mx40 mx246(.c0sm_b0m_v0m_n11(c0sm_b0m_v0m_n11), .c0sm_b0m_v0m_n262(c0sm_b0m_v0m_n262), .c0sm_b0m_v0m_n263(c0sm_b0m_v0m_n263), .clk(clk), .c0sm_b0m_rdata_0_(c0sm_b0m_rdata[0]), .c0sm_b0m_rdata_1_(c0sm_b0m_rdata[1]));
  /*CASIO@<instance>
     <id>mx247</id>
     <module>reg_mx41</module>
     <compmap>F1:c0nm_b0m_v0m_u67, F2:c0nm_b0m_v0m_u65, F3:c0nm_b0m_v0m_buffers1_reg_0_, F4:c0nm_b0m_v0m_buffers1_reg_1_, </compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  reg_mx41 mx247(.c0nm_b0m_v0m_n101(c0nm_b0m_v0m_n101), .c0nm_b0m_v0m_n97(c0nm_b0m_v0m_n97), .c0nm_b0m_v0m_n98(c0nm_b0m_v0m_n98), .clk(clk), .c0nm_b0m_v0m_n60(c0nm_b0m_v0m_n60), .c0nm_b0m_v0m_n61(c0nm_b0m_v0m_n61));
  /*CASIO@<instance>
     <id>mx248</id>
     <module>reg_mx42</module>
     <compmap>F1:c0sm_b0m_v0m_u67, F2:c0sm_b0m_v0m_u65, F3:c0sm_b0m_v0m_buffers1_reg_0_, F4:c0sm_b0m_v0m_buffers1_reg_1_, </compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  reg_mx42 mx248(.c0sm_b0m_v0m_n101(c0sm_b0m_v0m_n101), .c0sm_b0m_v0m_n97(c0sm_b0m_v0m_n97), .c0sm_b0m_v0m_n98(c0sm_b0m_v0m_n98), .clk(clk), .c0sm_b0m_v0m_n343(c0sm_b0m_v0m_n343), .c0sm_b0m_v0m_n344(c0sm_b0m_v0m_n344));
  /*CASIO@<instance>
     <id>mx249</id>
     <module>reg_mx43</module>
     <compmap>F1:c0nm_b0m_v0m_u207, F2:c0nm_b0m_v0m_u206, F3:c0nm_b0m_v0m_u205, F4:c0nm_b0m_v0m_u204, F5:c0nm_b0m_v0m_u203, F6:c0nm_b0m_v0m_u202, F7:c0nm_b0m_v0m_u201, F8:c0nm_b0m_v0m_u200, F9:c0nm_b0m_v0m_u199, F10:c0nm_b0m_v0m_u198, F11:c0nm_b0m_v0m_rdata_reg_10_, F12:c0nm_b0m_v0m_rdata_reg_11_, F13:c0nm_b0m_v0m_rdata_reg_2_, F14:c0nm_b0m_v0m_rdata_reg_3_, F15:c0nm_b0m_v0m_rdata_reg_4_, F16:c0nm_b0m_v0m_rdata_reg_5_, F17:c0nm_b0m_v0m_rdata_reg_6_, F18:c0nm_b0m_v0m_rdata_reg_7_, F19:c0nm_b0m_v0m_rdata_reg_8_, F20:c0nm_b0m_v0m_rdata_reg_9_, </compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  reg_mx43 mx249(.c0nm_b0m_headflit_10_(c0nm_b0m_headflit_10_), .c0nm_b0m_headflit_11_(c0nm_b0m_headflit_11_), .c0nm_b0m_headflit_8_(c0nm_b0m_headflit_8_), .c0nm_b0m_headflit_9_(c0nm_b0m_headflit_9_), .c0nm_b0m_v0m_n10(c0nm_b0m_v0m_n10), .c0nm_b0m_v0m_n11(c0nm_b0m_v0m_n11), .c0nm_headflit_2_(c0nm_headflit[2]), .c0nm_headflit_3_(c0nm_headflit[3]), .c0nm_headflit_4_(c0nm_headflit[4]), .c0nm_headflit_5_(c0nm_headflit[5]), .c0nm_headflit_6_(c0nm_headflit[6]), .c0nm_headflit_7_(c0nm_headflit[7]), .clk(clk), .c0nm_b0m_rdata_10_(c0nm_b0m_rdata[10]), .c0nm_b0m_rdata_11_(c0nm_b0m_rdata[11]), .c0nm_b0m_rdata_2_(c0nm_b0m_rdata[2]), .c0nm_b0m_rdata_3_(c0nm_b0m_rdata[3]), .c0nm_b0m_rdata_4_(c0nm_b0m_rdata[4]), .c0nm_b0m_rdata_5_(c0nm_b0m_rdata[5]), .c0nm_b0m_rdata_6_(c0nm_b0m_rdata[6]), .c0nm_b0m_rdata_7_(c0nm_b0m_rdata[7]), .c0nm_b0m_rdata_8_(c0nm_b0m_rdata[8]), .c0nm_b0m_rdata_9_(c0nm_b0m_rdata[9]));
  /*CASIO@<instance>
     <id>mx250</id>
     <module>reg_mx44</module>
     <compmap>F1:c0sm_b0m_v0m_u207, F2:c0sm_b0m_v0m_u206, F3:c0sm_b0m_v0m_u205, F4:c0sm_b0m_v0m_u204, F5:c0sm_b0m_v0m_u203, F6:c0sm_b0m_v0m_u202, F7:c0sm_b0m_v0m_u201, F8:c0sm_b0m_v0m_u200, F9:c0sm_b0m_v0m_u199, F10:c0sm_b0m_v0m_u198, F11:c0sm_b0m_v0m_rdata_reg_10_, F12:c0sm_b0m_v0m_rdata_reg_11_, F13:c0sm_b0m_v0m_rdata_reg_2_, F14:c0sm_b0m_v0m_rdata_reg_3_, F15:c0sm_b0m_v0m_rdata_reg_4_, F16:c0sm_b0m_v0m_rdata_reg_5_, F17:c0sm_b0m_v0m_rdata_reg_6_, F18:c0sm_b0m_v0m_rdata_reg_7_, F19:c0sm_b0m_v0m_rdata_reg_8_, F20:c0sm_b0m_v0m_rdata_reg_9_, </compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  reg_mx44 mx250(.c0sm_b0m_headflit_10_(c0sm_b0m_headflit_10_), .c0sm_b0m_headflit_11_(c0sm_b0m_headflit_11_), .c0sm_b0m_headflit_8_(c0sm_b0m_headflit_8_), .c0sm_b0m_headflit_9_(c0sm_b0m_headflit_9_), .c0sm_b0m_v0m_n10(c0sm_b0m_v0m_n10), .c0sm_b0m_v0m_n11(c0sm_b0m_v0m_n11), .c0sm_headflit_2_(c0sm_headflit[2]), .c0sm_headflit_3_(c0sm_headflit[3]), .c0sm_headflit_4_(c0sm_headflit[4]), .c0sm_headflit_5_(c0sm_headflit[5]), .c0sm_headflit_6_(c0sm_headflit[6]), .c0sm_headflit_7_(c0sm_headflit[7]), .clk(clk), .c0sm_b0m_rdata_10_(c0sm_b0m_rdata[10]), .c0sm_b0m_rdata_11_(c0sm_b0m_rdata[11]), .c0sm_b0m_rdata_2_(c0sm_b0m_rdata[2]), .c0sm_b0m_rdata_3_(c0sm_b0m_rdata[3]), .c0sm_b0m_rdata_4_(c0sm_b0m_rdata[4]), .c0sm_b0m_rdata_5_(c0sm_b0m_rdata[5]), .c0sm_b0m_rdata_6_(c0sm_b0m_rdata[6]), .c0sm_b0m_rdata_7_(c0sm_b0m_rdata[7]), .c0sm_b0m_rdata_8_(c0sm_b0m_rdata[8]), .c0sm_b0m_rdata_9_(c0sm_b0m_rdata[9]));
  /*CASIO@<instance>
     <id>mx251</id>
     <module>reg_mx45</module>
     <compmap>F1:c0nm_b0m_v0m_u78, F2:c0nm_b0m_v0m_u77, F3:c0nm_b0m_v0m_u76, F4:c0nm_b0m_v0m_u75, F5:c0nm_b0m_v0m_u74, F6:c0nm_b0m_v0m_u73, F7:c0nm_b0m_v0m_u72, F8:c0nm_b0m_v0m_u71, F9:c0nm_b0m_v0m_u70, F10:c0nm_b0m_v0m_u69, F11:c0nm_b0m_v0m_buffers1_reg_2_, F12:c0nm_b0m_v0m_buffers1_reg_3_, F13:c0nm_b0m_v0m_buffers1_reg_4_, F14:c0nm_b0m_v0m_buffers1_reg_5_, F15:c0nm_b0m_v0m_buffers1_reg_6_, F16:c0nm_b0m_v0m_buffers1_reg_7_, F17:c0nm_b0m_v0m_buffers1_reg_8_, F18:c0nm_b0m_v0m_buffers1_reg_9_, F19:c0nm_b0m_v0m_buffers1_reg_10_, F20:c0nm_b0m_v0m_buffers1_reg_11_, </compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  reg_mx45 mx251(.c0nm_b0m_v0m_n102(c0nm_b0m_v0m_n102), .c0nm_b0m_v0m_n103(c0nm_b0m_v0m_n103), .c0nm_b0m_v0m_n17(c0nm_b0m_v0m_n17), .c0nm_b0m_v0m_n19(c0nm_b0m_v0m_n19), .c0nm_b0m_v0m_n33(c0nm_b0m_v0m_n33), .c0nm_b0m_v0m_n34(c0nm_b0m_v0m_n34), .c0nm_b0m_v0m_n36(c0nm_b0m_v0m_n36), .c0nm_b0m_v0m_n37(c0nm_b0m_v0m_n37), .c0nm_b0m_v0m_n39(c0nm_b0m_v0m_n39), .c0nm_b0m_v0m_n40(c0nm_b0m_v0m_n40), .c0nm_b0m_v0m_n42(c0nm_b0m_v0m_n42), .c0nm_b0m_v0m_n43(c0nm_b0m_v0m_n43), .c0nm_b0m_v0m_n45(c0nm_b0m_v0m_n45), .c0nm_b0m_v0m_n46(c0nm_b0m_v0m_n46), .c0nm_b0m_v0m_n48(c0nm_b0m_v0m_n48), .c0nm_b0m_v0m_n49(c0nm_b0m_v0m_n49), .c0nm_b0m_v0m_n63(c0nm_b0m_v0m_n63), .c0nm_b0m_v0m_n64(c0nm_b0m_v0m_n64), .c0nm_b0m_v0m_n66(c0nm_b0m_v0m_n66), .c0nm_b0m_v0m_n67(c0nm_b0m_v0m_n67), .c0nm_b0m_v0m_n69(c0nm_b0m_v0m_n69), .c0nm_b0m_v0m_n70(c0nm_b0m_v0m_n70), .c0nm_b0m_v0m_n98(c0nm_b0m_v0m_n98), .clk(clk), .c0nm_b0m_v0m_n50(c0nm_b0m_v0m_n50), .c0nm_b0m_v0m_n51(c0nm_b0m_v0m_n51), .c0nm_b0m_v0m_n52(c0nm_b0m_v0m_n52), .c0nm_b0m_v0m_n53(c0nm_b0m_v0m_n53), .c0nm_b0m_v0m_n54(c0nm_b0m_v0m_n54), .c0nm_b0m_v0m_n55(c0nm_b0m_v0m_n55), .c0nm_b0m_v0m_n56(c0nm_b0m_v0m_n56), .c0nm_b0m_v0m_n57(c0nm_b0m_v0m_n57), .c0nm_b0m_v0m_n58(c0nm_b0m_v0m_n58), .c0nm_b0m_v0m_n59(c0nm_b0m_v0m_n59));
  /*CASIO@<instance>
     <id>mx252</id>
     <module>reg_mx46</module>
     <compmap>F1:c0sm_b0m_v0m_u78, F2:c0sm_b0m_v0m_u77, F3:c0sm_b0m_v0m_u76, F4:c0sm_b0m_v0m_u75, F5:c0sm_b0m_v0m_u74, F6:c0sm_b0m_v0m_u73, F7:c0sm_b0m_v0m_u72, F8:c0sm_b0m_v0m_u71, F9:c0sm_b0m_v0m_u70, F10:c0sm_b0m_v0m_u69, F11:c0sm_b0m_v0m_buffers1_reg_2_, F12:c0sm_b0m_v0m_buffers1_reg_3_, F13:c0sm_b0m_v0m_buffers1_reg_4_, F14:c0sm_b0m_v0m_buffers1_reg_5_, F15:c0sm_b0m_v0m_buffers1_reg_6_, F16:c0sm_b0m_v0m_buffers1_reg_7_, F17:c0sm_b0m_v0m_buffers1_reg_8_, F18:c0sm_b0m_v0m_buffers1_reg_9_, F19:c0sm_b0m_v0m_buffers1_reg_10_, F20:c0sm_b0m_v0m_buffers1_reg_11_, </compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  reg_mx46 mx252(.c0sm_b0m_v0m_n102(c0sm_b0m_v0m_n102), .c0sm_b0m_v0m_n103(c0sm_b0m_v0m_n103), .c0sm_b0m_v0m_n17(c0sm_b0m_v0m_n17), .c0sm_b0m_v0m_n19(c0sm_b0m_v0m_n19), .c0sm_b0m_v0m_n33(c0sm_b0m_v0m_n33), .c0sm_b0m_v0m_n34(c0sm_b0m_v0m_n34), .c0sm_b0m_v0m_n36(c0sm_b0m_v0m_n36), .c0sm_b0m_v0m_n37(c0sm_b0m_v0m_n37), .c0sm_b0m_v0m_n39(c0sm_b0m_v0m_n39), .c0sm_b0m_v0m_n40(c0sm_b0m_v0m_n40), .c0sm_b0m_v0m_n42(c0sm_b0m_v0m_n42), .c0sm_b0m_v0m_n43(c0sm_b0m_v0m_n43), .c0sm_b0m_v0m_n45(c0sm_b0m_v0m_n45), .c0sm_b0m_v0m_n46(c0sm_b0m_v0m_n46), .c0sm_b0m_v0m_n48(c0sm_b0m_v0m_n48), .c0sm_b0m_v0m_n49(c0sm_b0m_v0m_n49), .c0sm_b0m_v0m_n63(c0sm_b0m_v0m_n63), .c0sm_b0m_v0m_n64(c0sm_b0m_v0m_n64), .c0sm_b0m_v0m_n66(c0sm_b0m_v0m_n66), .c0sm_b0m_v0m_n67(c0sm_b0m_v0m_n67), .c0sm_b0m_v0m_n69(c0sm_b0m_v0m_n69), .c0sm_b0m_v0m_n70(c0sm_b0m_v0m_n70), .c0sm_b0m_v0m_n98(c0sm_b0m_v0m_n98), .clk(clk), .c0sm_b0m_v0m_n345(c0sm_b0m_v0m_n345), .c0sm_b0m_v0m_n346(c0sm_b0m_v0m_n346), .c0sm_b0m_v0m_n347(c0sm_b0m_v0m_n347), .c0sm_b0m_v0m_n348(c0sm_b0m_v0m_n348), .c0sm_b0m_v0m_n349(c0sm_b0m_v0m_n349), .c0sm_b0m_v0m_n350(c0sm_b0m_v0m_n350), .c0sm_b0m_v0m_n351(c0sm_b0m_v0m_n351), .c0sm_b0m_v0m_n352(c0sm_b0m_v0m_n352), .c0sm_b0m_v0m_n353(c0sm_b0m_v0m_n353), .c0sm_b0m_v0m_n354(c0sm_b0m_v0m_n354));
  /*CASIO@<instance>
     <id>mx259</id>
     <module>decoder24_mx47</module>
     <compmap>F1:d0m_u2, F2:d0m_u1</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  decoder24_mx47 mx259(.swalloc_resp_0_0_(swalloc_resp_0[0]), .swalloc_resp_1_0_(swalloc_resp_1[0]), .colsel0_0_(colsel0[0]), .colsel0_1_(colsel0[1]));
  /*CASIO@<instance>
     <id>mx260</id>
     <module>decoder24_mx48</module>
     <compmap>F1:d1m_u2, F2:d1m_u1</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  decoder24_mx48 mx260(.swalloc_resp_0_1_(swalloc_resp_0[1]), .swalloc_resp_1_1_(swalloc_resp_1[1]), .colsel1_0_(colsel1[0]), .colsel1_1_(colsel1[1]));
  /*CASIO@<instance>
     <id>mx261</id>
     <module>decoder24_mx49</module>
     <compmap>F1:s0m_o0nm_u29, F2:s0m_o0nm_u22</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  decoder24_mx49 mx261(.s0m_o0nm_state_credits_0_(s0m_o0nm_state_credits_0_), .s0m_o0nm_state_credits_1_(s0m_o0nm_state_credits_1_), .s0m_o0nm_n18(s0m_o0nm_n18), .s0m_o0nm_n22(s0m_o0nm_n22));
  /*CASIO@<instance>
     <id>mx262</id>
     <module>decoder24_mx50</module>
     <compmap>F1:s0m_o0sm_u29, F2:s0m_o0sm_u22</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  decoder24_mx50 mx262(.s0m_o0sm_state_credits_0_(s0m_o0sm_state_credits_0_), .s0m_o0sm_state_credits_1_(s0m_o0sm_state_credits_1_), .s0m_o0sm_n18(s0m_o0sm_n18), .s0m_o0sm_n22(s0m_o0sm_n22));
  /*CASIO@<instance>
     <id>mx271</id>
     <module>decoder38_mx51</module>
     <compmap>F1:s0m_o0nm_u27, F2:s0m_o0nm_u13, F3:s0m_o0nm_u12</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  decoder38_mx51 mx271(.creditin_0(creditin_0), .s0m_o0nm_n12(s0m_o0nm_n12), .s0m_o0nm_n9(s0m_o0nm_n9), .s0m_o0nm_n20(s0m_o0nm_n20), .s0m_o0nm_n6(s0m_o0nm_n6));
  /*CASIO@<instance>
     <id>mx272</id>
     <module>decoder38_mx52</module>
     <compmap>F1:s0m_o0sm_u27, F2:s0m_o0sm_u13, F3:s0m_o0sm_u12</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  decoder38_mx52 mx272(.creditin_1(creditin_1), .s0m_o0sm_n12(s0m_o0sm_n12), .s0m_o0sm_n9(s0m_o0sm_n9), .s0m_o0sm_n20(s0m_o0sm_n20), .s0m_o0sm_n6(s0m_o0sm_n6));
  /*CASIO@<instance>
     <id>mx276</id>
     <module>decoder38_mx53</module>
     <compmap>F1:c0nm_b0m_v0m_u193, F2:c0nm_b0m_v0m_u192, F3:c0nm_b0m_v0m_u189, F4:c0nm_b0m_v0m_u188, F5:c0nm_b0m_v0m_u186, F6:c0nm_b0m_v0m_u166, F7:c0nm_b0m_v0m_u165, F8:c0nm_b0m_v0m_u164, F9:c0nm_b0m_v0m_u80, F10:c0nm_b0m_v0m_u61</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  decoder38_mx53 mx276(.c0nm_b0m_v0m_n9(c0nm_b0m_v0m_n9), .c0nm_b0m_v0m_tail_0_(c0nm_b0m_v0m_tail_0_), .c0nm_b0m_v0m_tail_1_(c0nm_b0m_v0m_tail_1_), .c0nm_b0m_v0m_n100(c0nm_b0m_v0m_n100), .c0nm_b0m_v0m_n109(c0nm_b0m_v0m_n109), .c0nm_b0m_v0m_n78(c0nm_b0m_v0m_n78), .c0nm_b0m_v0m_n93(c0nm_b0m_v0m_n93), .c0nm_b0m_v0m_n94(c0nm_b0m_v0m_n94), .c0nm_b0m_v0m_n95(c0nm_b0m_v0m_n95));
  /*CASIO@<instance>
     <id>mx281</id>
     <module>decoder38_mx54</module>
     <compmap>F1:c0sm_b0m_v0m_u193, F2:c0sm_b0m_v0m_u192, F3:c0sm_b0m_v0m_u189, F4:c0sm_b0m_v0m_u188, F5:c0sm_b0m_v0m_u186, F6:c0sm_b0m_v0m_u166, F7:c0sm_b0m_v0m_u165, F8:c0sm_b0m_v0m_u164, F9:c0sm_b0m_v0m_u80, F10:c0sm_b0m_v0m_u61</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  decoder38_mx54 mx281(.c0sm_b0m_v0m_n355(c0sm_b0m_v0m_n355), .c0sm_b0m_v0m_tail_0_(c0sm_b0m_v0m_tail_0_), .c0sm_b0m_v0m_tail_1_(c0sm_b0m_v0m_tail_1_), .c0sm_b0m_v0m_n100(c0sm_b0m_v0m_n100), .c0sm_b0m_v0m_n109(c0sm_b0m_v0m_n109), .c0sm_b0m_v0m_n78(c0sm_b0m_v0m_n78), .c0sm_b0m_v0m_n93(c0sm_b0m_v0m_n93), .c0sm_b0m_v0m_n94(c0sm_b0m_v0m_n94), .c0sm_b0m_v0m_n95(c0sm_b0m_v0m_n95));
  /*CASIO@<instance>
     <id>mx309</id>
     <module>decoder416_mx55</module>
     <compmap>F1:c0nm_b0m_v0m_u278, F2:c0nm_b0m_v0m_u277, F3:c0nm_b0m_v0m_u276, F4:c0nm_b0m_v0m_u272, F5:c0nm_b0m_v0m_u271, F6:c0nm_b0m_v0m_u177, F7:c0nm_b0m_v0m_u176, F8:c0nm_b0m_v0m_u173, F9:c0nm_b0m_v0m_u172, F10:c0nm_b0m_v0m_u171</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  decoder416_mx55 mx309(.c0nm_b0m_v0m_head_0_(c0nm_b0m_v0m_head_0_), .c0nm_b0m_v0m_head_1_(c0nm_b0m_v0m_head_1_), .c0nm_b0m_v0m_head_2_(c0nm_b0m_v0m_head_2_), .debitout_0(debitout_0), .c0nm_b0m_v0m_n110(c0nm_b0m_v0m_n110), .c0nm_b0m_v0m_n113(c0nm_b0m_v0m_n113), .c0nm_b0m_v0m_n115(c0nm_b0m_v0m_n115));
  /*CASIO@<instance>
     <id>mx316</id>
     <module>decoder416_mx56</module>
     <compmap>F1:c0sm_b0m_v0m_u278, F2:c0sm_b0m_v0m_u277, F3:c0sm_b0m_v0m_u276, F4:c0sm_b0m_v0m_u272, F5:c0sm_b0m_v0m_u271, F6:c0sm_b0m_v0m_u177, F7:c0sm_b0m_v0m_u176, F8:c0sm_b0m_v0m_u173, F9:c0sm_b0m_v0m_u172, F10:c0sm_b0m_v0m_u171</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  decoder416_mx56 mx316(.c0sm_b0m_v0m_head_0_(c0sm_b0m_v0m_head_0_), .c0sm_b0m_v0m_head_1_(c0sm_b0m_v0m_head_1_), .c0sm_b0m_v0m_head_2_(c0sm_b0m_v0m_head_2_), .debitout_1(debitout_1), .c0sm_b0m_v0m_n110(c0sm_b0m_v0m_n110), .c0sm_b0m_v0m_n113(c0sm_b0m_v0m_n113), .c0sm_b0m_v0m_n115(c0sm_b0m_v0m_n115));
  /*CASIO@<instance>
     <id>mx319</id>
     <module>and2gate_mx57</module>
     <compmap>F1:c0nm_r0m_u16, F2:c0sm_r0m_u16</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  and2gate_mx57 mx319(.c0nm_r0m_n15(c0nm_r0m_n15), .c0sm_r0m_n15(c0sm_r0m_n15), .currx_1_(currx[1]), .c0nm_r0m_n16(c0nm_r0m_n16), .c0sm_r0m_n16(c0sm_r0m_n16));
  /*CASIO@<instance>
     <id>mx320</id>
     <module>and2gate_mx58</module>
     <compmap>F1:c0nm_b0m_u13, F2:c0nm_b0m_u12, F3:c0nm_b0m_u11, F4:c0nm_b0m_u10, F5:c0nm_b0m_u9, F6:c0nm_b0m_u8, F7:c0nm_b0m_u7, F8:c0nm_b0m_u6, F9:c0nm_b0m_u5, F10:c0nm_b0m_u4</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  and2gate_mx58 mx320(.c0nm_b0m_n1(c0nm_b0m_n1), .flitin_0_10_(flitin_0[10]), .flitin_0_11_(flitin_0[11]), .flitin_0_2_(flitin_0[2]), .flitin_0_3_(flitin_0[3]), .flitin_0_4_(flitin_0[4]), .flitin_0_5_(flitin_0[5]), .flitin_0_6_(flitin_0[6]), .flitin_0_7_(flitin_0[7]), .flitin_0_8_(flitin_0[8]), .flitin_0_9_(flitin_0[9]), .c0nm_b0m_wdata_10_(c0nm_b0m_wdata_10_), .c0nm_b0m_wdata_11_(c0nm_b0m_wdata_11_), .c0nm_b0m_wdata_2_(c0nm_b0m_wdata_2_), .c0nm_b0m_wdata_3_(c0nm_b0m_wdata_3_), .c0nm_b0m_wdata_4_(c0nm_b0m_wdata_4_), .c0nm_b0m_wdata_5_(c0nm_b0m_wdata_5_), .c0nm_b0m_wdata_6_(c0nm_b0m_wdata_6_), .c0nm_b0m_wdata_7_(c0nm_b0m_wdata_7_), .c0nm_b0m_wdata_8_(c0nm_b0m_wdata_8_), .c0nm_b0m_wdata_9_(c0nm_b0m_wdata_9_));
  /*CASIO@<instance>
     <id>mx321</id>
     <module>and2gate_mx59</module>
     <compmap>F1:c0nm_b0m_u25, F2:c0nm_b0m_u24, F3:c0nm_b0m_u22, F4:c0nm_b0m_u21, F5:c0nm_b0m_u20, F6:c0nm_b0m_u19, F7:c0nm_b0m_u18, F8:c0nm_b0m_u17, F9:c0nm_b0m_u16, F10:c0nm_b0m_u15</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  and2gate_mx59 mx321(.c0nm_b0m_dqenablereg(c0nm_b0m_dqenablereg), .c0nm_b0m_rdata_10_(c0nm_b0m_rdata[10]), .c0nm_b0m_rdata_11_(c0nm_b0m_rdata[11]), .c0nm_b0m_rdata_2_(c0nm_b0m_rdata[2]), .c0nm_b0m_rdata_3_(c0nm_b0m_rdata[3]), .c0nm_b0m_rdata_4_(c0nm_b0m_rdata[4]), .c0nm_b0m_rdata_5_(c0nm_b0m_rdata[5]), .c0nm_b0m_rdata_6_(c0nm_b0m_rdata[6]), .c0nm_b0m_rdata_7_(c0nm_b0m_rdata[7]), .c0nm_b0m_rdata_8_(c0nm_b0m_rdata[8]), .c0nm_b0m_rdata_9_(c0nm_b0m_rdata[9]), .flitout_switch_0_10_(flitout_switch_0[10]), .flitout_switch_0_11_(flitout_switch_0[11]), .flitout_switch_0_2_(flitout_switch_0[2]), .flitout_switch_0_3_(flitout_switch_0[3]), .flitout_switch_0_4_(flitout_switch_0[4]), .flitout_switch_0_5_(flitout_switch_0[5]), .flitout_switch_0_6_(flitout_switch_0[6]), .flitout_switch_0_7_(flitout_switch_0[7]), .flitout_switch_0_8_(flitout_switch_0[8]), .flitout_switch_0_9_(flitout_switch_0[9]));
  /*CASIO@<instance>
     <id>mx324</id>
     <module>and2gate_mx60</module>
     <compmap>F1:c0nm_v0m_u5, F2:s0m_u10</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  and2gate_mx60 mx324(.c0nm_v0m_n5(c0nm_v0m_n5), .s0m_elig_1_(s0m_elig_1_), .swalloc_req_0_1_(swalloc_req_0[1]), .c0nm_v0m_n3(c0nm_v0m_n3), .s0m_request0_1_(s0m_request0[1]));
  /*CASIO@<instance>
     <id>mx325</id>
     <module>and2gate_mx61</module>
     <compmap>F1:c0nm_v0m_u8, F2:s0m_u11</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  and2gate_mx61 mx325(.c0nm_v0m_n5(c0nm_v0m_n5), .s0m_elig_0_(s0m_elig_0_), .swalloc_req_0_0_(swalloc_req_0[0]), .c0nm_v0m_n7(c0nm_v0m_n7), .s0m_request0_0_(s0m_request0[0]));
  /*CASIO@<instance>
     <id>mx326</id>
     <module>and2gate_mx62</module>
     <compmap>F1:c0sm_b0m_u13, F2:c0sm_b0m_u12, F3:c0sm_b0m_u11, F4:c0sm_b0m_u10, F5:c0sm_b0m_u9, F6:c0sm_b0m_u8, F7:c0sm_b0m_u7, F8:c0sm_b0m_u6, F9:c0sm_b0m_u5, F10:c0sm_b0m_u4</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  and2gate_mx62 mx326(.c0sm_b0m_n2(c0sm_b0m_n2), .flitin_1_10_(flitin_1[10]), .flitin_1_11_(flitin_1[11]), .flitin_1_2_(flitin_1[2]), .flitin_1_3_(flitin_1[3]), .flitin_1_4_(flitin_1[4]), .flitin_1_5_(flitin_1[5]), .flitin_1_6_(flitin_1[6]), .flitin_1_7_(flitin_1[7]), .flitin_1_8_(flitin_1[8]), .flitin_1_9_(flitin_1[9]), .c0sm_b0m_wdata_10_(c0sm_b0m_wdata_10_), .c0sm_b0m_wdata_11_(c0sm_b0m_wdata_11_), .c0sm_b0m_wdata_2_(c0sm_b0m_wdata_2_), .c0sm_b0m_wdata_3_(c0sm_b0m_wdata_3_), .c0sm_b0m_wdata_4_(c0sm_b0m_wdata_4_), .c0sm_b0m_wdata_5_(c0sm_b0m_wdata_5_), .c0sm_b0m_wdata_6_(c0sm_b0m_wdata_6_), .c0sm_b0m_wdata_7_(c0sm_b0m_wdata_7_), .c0sm_b0m_wdata_8_(c0sm_b0m_wdata_8_), .c0sm_b0m_wdata_9_(c0sm_b0m_wdata_9_));
  /*CASIO@<instance>
     <id>mx327</id>
     <module>and2gate_mx63</module>
     <compmap>F1:c0sm_b0m_u25, F2:c0sm_b0m_u24, F3:c0sm_b0m_u22, F4:c0sm_b0m_u21, F5:c0sm_b0m_u20, F6:c0sm_b0m_u19, F7:c0sm_b0m_u18, F8:c0sm_b0m_u17, F9:c0sm_b0m_u16, F10:c0sm_b0m_u15</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  and2gate_mx63 mx327(.c0sm_b0m_dqenablereg(c0sm_b0m_dqenablereg), .c0sm_b0m_rdata_10_(c0sm_b0m_rdata[10]), .c0sm_b0m_rdata_11_(c0sm_b0m_rdata[11]), .c0sm_b0m_rdata_2_(c0sm_b0m_rdata[2]), .c0sm_b0m_rdata_3_(c0sm_b0m_rdata[3]), .c0sm_b0m_rdata_4_(c0sm_b0m_rdata[4]), .c0sm_b0m_rdata_5_(c0sm_b0m_rdata[5]), .c0sm_b0m_rdata_6_(c0sm_b0m_rdata[6]), .c0sm_b0m_rdata_7_(c0sm_b0m_rdata[7]), .c0sm_b0m_rdata_8_(c0sm_b0m_rdata[8]), .c0sm_b0m_rdata_9_(c0sm_b0m_rdata[9]), .flitout_switch_1_10_(flitout_switch_1[10]), .flitout_switch_1_11_(flitout_switch_1[11]), .flitout_switch_1_2_(flitout_switch_1[2]), .flitout_switch_1_3_(flitout_switch_1[3]), .flitout_switch_1_4_(flitout_switch_1[4]), .flitout_switch_1_5_(flitout_switch_1[5]), .flitout_switch_1_6_(flitout_switch_1[6]), .flitout_switch_1_7_(flitout_switch_1[7]), .flitout_switch_1_8_(flitout_switch_1[8]), .flitout_switch_1_9_(flitout_switch_1[9]));
  /*CASIO@<instance>
     <id>mx330</id>
     <module>and2gate_mx64</module>
     <compmap>F1:c0sm_v0m_u5, F2:s0m_u8</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  and2gate_mx64 mx330(.c0sm_v0m_n5(c0sm_v0m_n5), .s0m_elig_1_(s0m_elig_1_), .swalloc_req_1_1_(swalloc_req_1[1]), .c0sm_v0m_n3(c0sm_v0m_n3), .s0m_request1_1_(s0m_request1[1]));
  /*CASIO@<instance>
     <id>mx331</id>
     <module>and2gate_mx65</module>
     <compmap>F1:c0sm_v0m_u8, F2:s0m_u9</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  and2gate_mx65 mx331(.c0sm_v0m_n5(c0sm_v0m_n5), .s0m_elig_0_(s0m_elig_0_), .swalloc_req_1_0_(swalloc_req_1[0]), .c0sm_v0m_n7(c0sm_v0m_n7), .s0m_request1_0_(s0m_request1[0]));
  /*CASIO@<instance>
     <id>mx334</id>
     <module>or2gate_mx66</module>
     <compmap>F1:c0nm_r0m_u18, F2:c0sm_r0m_u18</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  or2gate_mx66 mx334(.c0nm_r0m_n9(c0nm_r0m_n9), .c0sm_r0m_n9(c0sm_r0m_n9), .currx_0_(currx[0]), .c0nm_r0m_n15(c0nm_r0m_n15), .c0sm_r0m_n15(c0sm_r0m_n15));
  /*CASIO@<instance>
     <id>mx335</id>
     <module>or2gate_mx67</module>
     <compmap>F1:c0nm_b0m_v0m_u262, F2:c0nm_b0m_v0m_u261, F3:c0nm_b0m_v0m_u197, F4:c0nm_b0m_v0m_u195, F5:c0nm_b0m_v0m_u179, F6:c0nm_b0m_v0m_u178, F7:c0nm_b0m_v0m_u83, F8:c0nm_b0m_v0m_u82, F9:c0nm_b0m_v0m_u64, F10:c0nm_b0m_v0m_u63, F11:c0nm_b0m_v0m_u7, F12:c0nm_b0m_v0m_u4, F13:c0nm_v0m_u38, F14:c0nm_v0m_u9, F15:c0sm_b0m_v0m_u262, F16:c0sm_b0m_v0m_u197, F17:c0sm_b0m_v0m_u195, F18:c0sm_b0m_v0m_u179, F19:c0sm_b0m_v0m_u178, F20:c0sm_b0m_v0m_u83, F21:c0sm_b0m_v0m_u82, F22:c0sm_b0m_v0m_u64, F23:c0sm_b0m_v0m_u63, F24:c0sm_b0m_v0m_u7, F25:c0sm_b0m_v0m_u4, F26:c0sm_v0m_u38, F27:c0sm_v0m_u9, F28:x0m_u8, F29:x0m_u7, F30:x0m_u6, F31:x0m_u5</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  or2gate_mx67 mx335(.c0nm_b0m_n1(c0nm_b0m_n1), .c0nm_b0m_v0m_n8(c0nm_b0m_v0m_n8), .c0nm_b0m_v0m_n93(c0nm_b0m_v0m_n93), .c0nm_b0m_v0m_n94(c0nm_b0m_v0m_n94), .c0nm_b0m_v0m_n95(c0nm_b0m_v0m_n95), .c0nm_headflit_0_(c0nm_headflit[0]), .c0nm_headflit_1_(c0nm_headflit[1]), .c0sm_b0m_n2(c0sm_b0m_n2), .c0sm_b0m_v0m_n8(c0sm_b0m_v0m_n8), .c0sm_b0m_v0m_n93(c0sm_b0m_v0m_n93), .c0sm_b0m_v0m_n94(c0sm_b0m_v0m_n94), .c0sm_b0m_v0m_n95(c0sm_b0m_v0m_n95), .c0sm_headflit_0_(c0sm_headflit[0]), .c0sm_headflit_1_(c0sm_headflit[1]), .colsel0_0_(colsel0[0]), .colsel0_1_(colsel0[1]), .colsel1_0_(colsel1[0]), .colsel1_1_(colsel1[1]), .reset(reset), .tailout_0(tailout_0), .tailout_1(tailout_1), .c0nm_b0m_v0m_n1(c0nm_b0m_v0m_n1), .c0nm_b0m_v0m_n102(c0nm_b0m_v0m_n102), .c0nm_b0m_v0m_n129(c0nm_b0m_v0m_n129), .c0nm_b0m_v0m_n2(c0nm_b0m_v0m_n2), .c0nm_b0m_v0m_n262(c0nm_b0m_v0m_n262), .c0nm_b0m_v0m_n263(c0nm_b0m_v0m_n263), .c0nm_b0m_v0m_n81(c0nm_b0m_v0m_n81), .c0nm_v0m_n1(c0nm_v0m_n1), .c0sm_b0m_v0m_n1(c0sm_b0m_v0m_n1), .c0sm_b0m_v0m_n102(c0sm_b0m_v0m_n102), .c0sm_b0m_v0m_n129(c0sm_b0m_v0m_n129), .c0sm_b0m_v0m_n2(c0sm_b0m_v0m_n2), .c0sm_b0m_v0m_n262(c0sm_b0m_v0m_n262), .c0sm_b0m_v0m_n263(c0sm_b0m_v0m_n263), .c0sm_b0m_v0m_n81(c0sm_b0m_v0m_n81), .c0sm_v0m_n1(c0sm_v0m_n1), .x0m_n3(x0m_n3), .x0m_n4(x0m_n4), .x0m_n5(x0m_n5), .x0m_n6(x0m_n6));
  /*CASIO@<instance>
     <id>mx336</id>
     <module>or2gate_mx68</module>
     <compmap>F1:c0nm_b0m_v0m_u191, F2:c0nm_b0m_v0m_u190, F3:c0nm_b0m_v0m_u182, F4:c0nm_b0m_v0m_u98</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  or2gate_mx68 mx336(.c0nm_b0m_n1(c0nm_b0m_n1), .c0nm_b0m_v0m_n28(c0nm_b0m_v0m_n28), .c0nm_b0m_v0m_n93(c0nm_b0m_v0m_n93), .c0nm_b0m_v0m_n116(c0nm_b0m_v0m_n116), .c0nm_b0m_v0m_n135(c0nm_b0m_v0m_n135));
  /*CASIO@<instance>
     <id>mx338</id>
     <module>or2gate_mx69</module>
     <compmap>F1:c0sm_b0m_v0m_u191, F2:c0sm_b0m_v0m_u190, F3:c0sm_b0m_v0m_u182, F4:c0sm_b0m_v0m_u98</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  or2gate_mx69 mx338(.c0sm_b0m_n2(c0sm_b0m_n2), .c0sm_b0m_v0m_n28(c0sm_b0m_v0m_n28), .c0sm_b0m_v0m_n93(c0sm_b0m_v0m_n93), .c0sm_b0m_v0m_n116(c0sm_b0m_v0m_n116), .c0sm_b0m_v0m_n135(c0sm_b0m_v0m_n135));
  /*CASIO@<instance>
     <id>mx341</id>
     <module>or2gate_mx70</module>
     <compmap>F1:x0m_u4, F2:x0m_bx0m_m1m_m4m_u1, F3:x0m_bx1m_m1m_m4m_u1</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  or2gate_mx70 mx341(.x0m_bx0m_m1m_int01(x0m_bx0m_m1m_int01), .x0m_bx1m_m1m_int01(x0m_bx1m_m1m_int01), .x0m_colsel1reg_1_(x0m_colsel1reg_1_), .flitout_1_0_(flitout_1[0]), .flitout_1_1_(flitout_1[1]));
  /*CASIO@<instance>
     <id>mx343</id>
     <module>nand2gate_mx71</module>
     <compmap>F1:c0nm_u3, F2:c0nm_b0m_u14</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  nand2gate_mx71 mx343(.flitin_0_0_(flitin_0[0]), .flitin_0_1_(flitin_0[1]), .c0nm_b0m_n1(c0nm_b0m_n1), .c0nm_n2(c0nm_n2));
  /*CASIO@<instance>
     <id>mx345</id>
     <module>nand2gate_mx72</module>
     <compmap>F1:c0sm_u3, F2:c0sm_b0m_u14</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  nand2gate_mx72 mx345(.flitin_1_0_(flitin_1[0]), .flitin_1_1_(flitin_1[1]), .c0sm_b0m_n2(c0sm_b0m_n2), .c0sm_n3(c0sm_n3));
  /*CASIO@<instance>
     <id>mx346</id>
     <module>nand2gate_mx73</module>
     <compmap>F1:c0nm_b0m_v0m_u31, F2:c0sm_b0m_v0m_u31, F3:s0m_o0nm_u23, F4:s0m_o0sm_u23</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  nand2gate_mx73 mx346(.c0nm_b0m_v0m_n26(c0nm_b0m_v0m_n26), .c0nm_b0m_v0m_n4(c0nm_b0m_v0m_n4), .c0sm_b0m_v0m_n26(c0sm_b0m_v0m_n26), .s0m_o0nm_n24(s0m_o0nm_n24), .s0m_o0sm_n24(s0m_o0sm_n24), .c0nm_b0m_v0m_n20(c0nm_b0m_v0m_n20), .c0sm_b0m_v0m_n20(c0sm_b0m_v0m_n20), .s0m_o0nm_n36(s0m_o0nm_n36), .s0m_o0sm_n36(s0m_o0sm_n36));
  /*CASIO@<instance>
     <id>mx347</id>
     <module>nand2gate_mx74</module>
     <compmap>F1:s0m_u7, F2:s0m_u4</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  nand2gate_mx74 mx347(.s0m_state_invc0_1_(s0m_state_invc0_1_), .s0m_state_invc1_1_(s0m_state_invc1_1_), .tailout_1(tailout_1), .s0m_n1(s0m_n1), .s0m_n3(s0m_n3));
  /*CASIO@<instance>
     <id>mx348</id>
     <module>nand2gate_mx75</module>
     <compmap>F1:s0m_u38, F2:s0m_u35</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  nand2gate_mx75 mx348(.debitout_1(debitout_1), .s0m_state_invc0_1_(s0m_state_invc0_1_), .s0m_state_invc1_1_(s0m_state_invc1_1_), .s0m_n20(s0m_n20), .s0m_n26(s0m_n26));
  /*CASIO@<instance>
     <id>mx349</id>
     <module>nand2gate_mx76</module>
     <compmap>F1:s0m_u31, F2:s0m_u26</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  nand2gate_mx76 mx349(.s0m_n16(s0m_n16), .s0m_outb0_1_(s0m_outb0_1_), .s0m_outb1_1_(s0m_outb1_1_), .s0m_n14(s0m_n14), .s0m_n18(s0m_n18));
  /*CASIO@<instance>
     <id>mx350</id>
     <module>nand2gate_mx77</module>
     <compmap>F1:s0m_u22, F2:s0m_u17</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  nand2gate_mx77 mx350(.s0m_n9(s0m_n9), .s0m_outb0_0_(s0m_outb0_0_), .s0m_outb1_0_(s0m_outb1_0_), .s0m_n11(s0m_n11), .s0m_n7(s0m_n7));
  /*CASIO@<instance>
     <id>mx353</id>
     <module>nor2gate_mx78</module>
     <compmap>F1:c0nm_u5, F2:c0nm_b0m_v0m_u209, F3:c0nm_b0m_v0m_u208, F4:c0nm_b0m_v0m_u10, F5:c0nm_v0m_u23, F6:c0nm_v0m_u17, F7:c0nm_v0m_u11, F8:c0sm_u5, F9:c0sm_b0m_v0m_u209, F10:c0sm_b0m_v0m_u208, F11:c0sm_b0m_v0m_u10, F12:c0sm_v0m_u23, F13:c0sm_v0m_u17, F14:c0sm_v0m_u11, F15:s0m_u32, F16:s0m_u23, F17:s0m_m0m_u4, F18:s0m_m1m_u4, F19:s0m_o0nm_u35, F20:s0m_o0nm_u14, F21:s0m_o0sm_u35, F22:s0m_o0sm_u14</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  nor2gate_mx78 mx353(.c0nm_b0m_n1(c0nm_b0m_n1), .c0nm_v0m_n10(c0nm_v0m_n10), .c0nm_v0m_n19(c0nm_v0m_n19), .c0nm_v0m_n27(c0nm_v0m_n27), .c0sm_b0m_n2(c0sm_b0m_n2), .c0sm_v0m_n10(c0sm_v0m_n10), .c0sm_v0m_n19(c0sm_v0m_n19), .c0sm_v0m_n27(c0sm_v0m_n27), .debitout_0(debitout_0), .debitout_1(debitout_1), .reset(reset), .s0m_m0m_n2(s0m_m0m_n2), .s0m_m1m_n2(s0m_m1m_n2), .s0m_o0nm_n13(s0m_o0nm_n13), .s0m_o0sm_n13(s0m_o0sm_n13), .s0m_tail_outvc0(s0m_tail_outvc0), .s0m_tail_outvc1(s0m_tail_outvc1), .tailout_0(tailout_0), .tailout_1(tailout_1), .c0nm_b0m_v0m_n10(c0nm_b0m_v0m_n10), .c0nm_b0m_v0m_n11(c0nm_b0m_v0m_n11), .c0nm_b0m_v0m_n8(c0nm_b0m_v0m_n8), .c0nm_v0m_n61(c0nm_v0m_n61), .c0nm_v0m_n62(c0nm_v0m_n62), .c0nm_v0m_n64(c0nm_v0m_n64), .c0sm_b0m_v0m_n10(c0sm_b0m_v0m_n10), .c0sm_b0m_v0m_n11(c0sm_b0m_v0m_n11), .c0sm_b0m_v0m_n8(c0sm_b0m_v0m_n8), .c0sm_v0m_n61(c0sm_v0m_n61), .c0sm_v0m_n62(c0sm_v0m_n62), .c0sm_v0m_n64(c0sm_v0m_n64), .creditout_0(creditout_0), .creditout_1(creditout_1), .s0m_m0m_n10(s0m_m0m_n10), .s0m_m1m_n10(s0m_m1m_n10), .s0m_n16(s0m_n16), .s0m_n9(s0m_n9), .s0m_o0nm_n3(s0m_o0nm_n3), .s0m_o0nm_n38(s0m_o0nm_n38), .s0m_o0sm_n3(s0m_o0sm_n3), .s0m_o0sm_n38(s0m_o0sm_n38));
  /*CASIO@<instance>
     <id>mx354</id>
     <module>nor2gate_mx79</module>
     <compmap>F1:c0nm_b0m_v0m_u187, F2:c0nm_b0m_v0m_u185</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  nor2gate_mx79 mx354(.c0nm_b0m_n1(c0nm_b0m_n1), .c0nm_b0m_v0m_n94(c0nm_b0m_v0m_n94), .c0nm_b0m_v0m_n95(c0nm_b0m_v0m_n95), .c0nm_b0m_v0m_n120(c0nm_b0m_v0m_n120), .c0nm_b0m_v0m_n121(c0nm_b0m_v0m_n121));
  /*CASIO@<instance>
     <id>mx356</id>
     <module>nor2gate_mx80</module>
     <compmap>F1:c0nm_b0m_u27, F2:c0nm_v0m_u30, F3:c0nm_v0m_u10</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  nor2gate_mx80 mx356(.c0nm_n2(c0nm_n2), .c0nm_v0m_n9(c0nm_v0m_n9), .reset(reset), .c0nm_b0m_n9(c0nm_b0m_n9), .c0nm_v0m_n13(c0nm_v0m_n13));
  /*CASIO@<instance>
     <id>mx358</id>
     <module>nor2gate_mx81</module>
     <compmap>F1:c0nm_v0m_u6, F2:c0nm_v0m_u3</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  nor2gate_mx81 mx358(.c0nm_v0m_n1(c0nm_v0m_n1), .c0nm_v0m_n2(c0nm_v0m_n2), .c0nm_v0m_n6(c0nm_v0m_n6), .c0nm_v0m_n30(c0nm_v0m_n30), .c0nm_v0m_n31(c0nm_v0m_n31));
  /*CASIO@<instance>
     <id>mx359</id>
     <module>nor2gate_mx82</module>
     <compmap>F1:c0sm_b0m_v0m_u187, F2:c0sm_b0m_v0m_u185</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  nor2gate_mx82 mx359(.c0sm_b0m_n2(c0sm_b0m_n2), .c0sm_b0m_v0m_n94(c0sm_b0m_v0m_n94), .c0sm_b0m_v0m_n95(c0sm_b0m_v0m_n95), .c0sm_b0m_v0m_n120(c0sm_b0m_v0m_n120), .c0sm_b0m_v0m_n121(c0sm_b0m_v0m_n121));
  /*CASIO@<instance>
     <id>mx361</id>
     <module>nor2gate_mx83</module>
     <compmap>F1:c0sm_b0m_u27, F2:c0sm_v0m_u30, F3:c0sm_v0m_u10</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  nor2gate_mx83 mx361(.c0sm_n3(c0sm_n3), .c0sm_v0m_n9(c0sm_v0m_n9), .reset(reset), .c0sm_b0m_n9(c0sm_b0m_n9), .c0sm_v0m_n13(c0sm_v0m_n13));
  /*CASIO@<instance>
     <id>mx363</id>
     <module>nor2gate_mx84</module>
     <compmap>F1:c0sm_v0m_u6, F2:c0sm_v0m_u3</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  nor2gate_mx84 mx363(.c0sm_v0m_n1(c0sm_v0m_n1), .c0sm_v0m_n2(c0sm_v0m_n2), .c0sm_v0m_n6(c0sm_v0m_n6), .c0sm_v0m_n32(c0sm_v0m_n32), .c0sm_v0m_n33(c0sm_v0m_n33));
  /*CASIO@<instance>
     <id>mx366</id>
     <module>mux_merged_mx85</module>
     <compmap>F1:c0nm_b0m_v0m_u92, F2:c0nm_b0m_v0m_u91, F3:c0nm_b0m_v0m_u85, F4:c0nm_b0m_v0m_u84</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux_merged_mx85 mx366(.c0nm_b0m_v0m_n105(c0nm_b0m_v0m_n105), .c0nm_b0m_v0m_n107(c0nm_b0m_v0m_n107), .c0nm_b0m_v0m_n108(c0nm_b0m_v0m_n108), .c0nm_b0m_v0m_n109(c0nm_b0m_v0m_n109), .c0nm_b0m_v0m_n122(c0nm_b0m_v0m_n122), .c0nm_b0m_v0m_n25(c0nm_b0m_v0m_n25), .c0nm_b0m_v0m_n27(c0nm_b0m_v0m_n27), .c0nm_b0m_v0m_n31(c0nm_b0m_v0m_n31), .c0nm_b0m_v0m_n32(c0nm_b0m_v0m_n32), .reset(reset), .c0nm_b0m_v0m_n218(c0nm_b0m_v0m_n218), .c0nm_b0m_v0m_n219(c0nm_b0m_v0m_n219));
  /*CASIO@<instance>
     <id>mx368</id>
     <module>mux_merged_mx86</module>
     <compmap>F1:c0nm_b0m_v0m_u38, F2:c0nm_b0m_v0m_u37, F3:c0nm_b0m_v0m_u35, F4:c0nm_b0m_v0m_u34</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux_merged_mx86 mx368(.c0nm_b0m_v0m_n25(c0nm_b0m_v0m_n25), .c0nm_b0m_v0m_n27(c0nm_b0m_v0m_n27), .c0nm_b0m_v0m_n31(c0nm_b0m_v0m_n31), .c0nm_b0m_v0m_n32(c0nm_b0m_v0m_n32), .c0nm_b0m_v0m_n74(c0nm_b0m_v0m_n74), .c0nm_b0m_v0m_n76(c0nm_b0m_v0m_n76), .c0nm_b0m_v0m_n77(c0nm_b0m_v0m_n77), .c0nm_b0m_v0m_n78(c0nm_b0m_v0m_n78), .c0nm_b0m_v0m_n79(c0nm_b0m_v0m_n79), .reset(reset), .c0nm_b0m_v0m_n242(c0nm_b0m_v0m_n242), .c0nm_b0m_v0m_n243(c0nm_b0m_v0m_n243));
  /*CASIO@<instance>
     <id>mx369</id>
     <module>mux_merged_mx87</module>
     <compmap>F1:c0nm_b0m_v0m_u21, F2:c0nm_b0m_v0m_u20, F3:c0nm_b0m_v0m_u19, F4:c0nm_b0m_v0m_u18</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux_merged_mx87 mx369(.c0nm_b0m_v0m_n22(c0nm_b0m_v0m_n22), .c0nm_b0m_v0m_n23(c0nm_b0m_v0m_n23), .c0nm_b0m_v0m_n25(c0nm_b0m_v0m_n25), .c0nm_b0m_v0m_n26(c0nm_b0m_v0m_n26), .c0nm_b0m_v0m_n27(c0nm_b0m_v0m_n27), .c0nm_b0m_v0m_n28(c0nm_b0m_v0m_n28), .c0nm_b0m_v0m_n29(c0nm_b0m_v0m_n29), .c0nm_b0m_v0m_n31(c0nm_b0m_v0m_n31), .c0nm_b0m_v0m_n32(c0nm_b0m_v0m_n32), .reset(reset), .c0nm_b0m_v0m_n253(c0nm_b0m_v0m_n253), .c0nm_b0m_v0m_n254(c0nm_b0m_v0m_n254));
  /*CASIO@<instance>
     <id>mx370</id>
     <module>mux_merged_mx88</module>
     <compmap>F1:c0sm_b0m_v0m_u92, F2:c0sm_b0m_v0m_u91, F3:c0sm_b0m_v0m_u85, F4:c0sm_b0m_v0m_u84</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux_merged_mx88 mx370(.c0sm_b0m_v0m_n105(c0sm_b0m_v0m_n105), .c0sm_b0m_v0m_n107(c0sm_b0m_v0m_n107), .c0sm_b0m_v0m_n108(c0sm_b0m_v0m_n108), .c0sm_b0m_v0m_n109(c0sm_b0m_v0m_n109), .c0sm_b0m_v0m_n122(c0sm_b0m_v0m_n122), .c0sm_b0m_v0m_n25(c0sm_b0m_v0m_n25), .c0sm_b0m_v0m_n27(c0sm_b0m_v0m_n27), .c0sm_b0m_v0m_n31(c0sm_b0m_v0m_n31), .c0sm_b0m_v0m_n32(c0sm_b0m_v0m_n32), .reset(reset), .c0sm_b0m_v0m_n319(c0sm_b0m_v0m_n319), .c0sm_b0m_v0m_n320(c0sm_b0m_v0m_n320));
  /*CASIO@<instance>
     <id>mx372</id>
     <module>mux_merged_mx89</module>
     <compmap>F1:c0sm_b0m_v0m_u38, F2:c0sm_b0m_v0m_u37, F3:c0sm_b0m_v0m_u35, F4:c0sm_b0m_v0m_u34</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux_merged_mx89 mx372(.c0sm_b0m_v0m_n25(c0sm_b0m_v0m_n25), .c0sm_b0m_v0m_n27(c0sm_b0m_v0m_n27), .c0sm_b0m_v0m_n31(c0sm_b0m_v0m_n31), .c0sm_b0m_v0m_n32(c0sm_b0m_v0m_n32), .c0sm_b0m_v0m_n74(c0sm_b0m_v0m_n74), .c0sm_b0m_v0m_n76(c0sm_b0m_v0m_n76), .c0sm_b0m_v0m_n77(c0sm_b0m_v0m_n77), .c0sm_b0m_v0m_n78(c0sm_b0m_v0m_n78), .c0sm_b0m_v0m_n79(c0sm_b0m_v0m_n79), .reset(reset), .c0sm_b0m_v0m_n295(c0sm_b0m_v0m_n295), .c0sm_b0m_v0m_n296(c0sm_b0m_v0m_n296));
  /*CASIO@<instance>
     <id>mx373</id>
     <module>mux_merged_mx90</module>
     <compmap>F1:c0sm_b0m_v0m_u21, F2:c0sm_b0m_v0m_u20, F3:c0sm_b0m_v0m_u19, F4:c0sm_b0m_v0m_u18</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux_merged_mx90 mx373(.c0sm_b0m_v0m_n22(c0sm_b0m_v0m_n22), .c0sm_b0m_v0m_n23(c0sm_b0m_v0m_n23), .c0sm_b0m_v0m_n25(c0sm_b0m_v0m_n25), .c0sm_b0m_v0m_n26(c0sm_b0m_v0m_n26), .c0sm_b0m_v0m_n27(c0sm_b0m_v0m_n27), .c0sm_b0m_v0m_n28(c0sm_b0m_v0m_n28), .c0sm_b0m_v0m_n29(c0sm_b0m_v0m_n29), .c0sm_b0m_v0m_n31(c0sm_b0m_v0m_n31), .c0sm_b0m_v0m_n32(c0sm_b0m_v0m_n32), .reset(reset), .c0sm_b0m_v0m_n284(c0sm_b0m_v0m_n284), .c0sm_b0m_v0m_n285(c0sm_b0m_v0m_n285));
  /*CASIO@<instance>
     <id>mx374</id>
     <module>mux_merged_mx91</module>
     <compmap>F1:c0nm_b0m_v0m_u256, F2:c0nm_b0m_v0m_u255, F3:c0nm_b0m_v0m_u251, F4:c0nm_b0m_v0m_u250, F5:c0nm_b0m_v0m_u246, F6:c0nm_b0m_v0m_u245, F7:c0nm_b0m_v0m_u236, F8:c0nm_b0m_v0m_u235, F9:c0nm_b0m_v0m_u221, F10:c0nm_b0m_v0m_u220, F11:c0nm_b0m_v0m_u216, F12:c0nm_b0m_v0m_u215, F13:c0nm_b0m_v0m_u211, F14:c0nm_b0m_v0m_u210</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux_merged_mx91 mx374(.c0nm_b0m_v0m_buffers0_10_(c0nm_b0m_v0m_buffers0_10_), .c0nm_b0m_v0m_buffers0_11_(c0nm_b0m_v0m_buffers0_11_), .c0nm_b0m_v0m_buffers0_2_(c0nm_b0m_v0m_buffers0_2_), .c0nm_b0m_v0m_buffers0_4_(c0nm_b0m_v0m_buffers0_4_), .c0nm_b0m_v0m_buffers0_7_(c0nm_b0m_v0m_buffers0_7_), .c0nm_b0m_v0m_buffers0_8_(c0nm_b0m_v0m_buffers0_8_), .c0nm_b0m_v0m_buffers0_9_(c0nm_b0m_v0m_buffers0_9_), .c0nm_b0m_v0m_n131(c0nm_b0m_v0m_n131), .c0nm_b0m_v0m_n134(c0nm_b0m_v0m_n134), .c0nm_b0m_v0m_n144(c0nm_b0m_v0m_n144), .c0nm_b0m_v0m_n147(c0nm_b0m_v0m_n147), .c0nm_b0m_v0m_n162(c0nm_b0m_v0m_n162), .c0nm_b0m_v0m_n165(c0nm_b0m_v0m_n165), .c0nm_b0m_v0m_n168(c0nm_b0m_v0m_n168), .c0nm_b0m_v0m_n171(c0nm_b0m_v0m_n171), .c0nm_b0m_v0m_n174(c0nm_b0m_v0m_n174), .c0nm_b0m_v0m_n177(c0nm_b0m_v0m_n177), .c0nm_b0m_v0m_n180(c0nm_b0m_v0m_n180), .c0nm_b0m_v0m_n183(c0nm_b0m_v0m_n183), .c0nm_b0m_v0m_n186(c0nm_b0m_v0m_n186), .c0nm_b0m_v0m_n187(c0nm_b0m_v0m_n187), .c0nm_b0m_v0m_n190(c0nm_b0m_v0m_n190), .c0nm_b0m_v0m_n192(c0nm_b0m_v0m_n192), .c0nm_b0m_v0m_n193(c0nm_b0m_v0m_n193), .c0nm_b0m_v0m_n21(c0nm_b0m_v0m_n21), .c0nm_b0m_v0m_n35(c0nm_b0m_v0m_n35), .c0nm_b0m_v0m_n41(c0nm_b0m_v0m_n41), .c0nm_b0m_v0m_n62(c0nm_b0m_v0m_n62), .c0nm_b0m_v0m_n65(c0nm_b0m_v0m_n65), .c0nm_b0m_v0m_n68(c0nm_b0m_v0m_n68), .c0nm_b0m_v0m_n71(c0nm_b0m_v0m_n71), .c0nm_b0m_v0m_n73(c0nm_b0m_v0m_n73), .c0nm_b0m_headflit_10_(c0nm_b0m_headflit_10_), .c0nm_b0m_headflit_11_(c0nm_b0m_headflit_11_), .c0nm_b0m_headflit_8_(c0nm_b0m_headflit_8_), .c0nm_b0m_headflit_9_(c0nm_b0m_headflit_9_), .c0nm_headflit_2_(c0nm_headflit[2]), .c0nm_headflit_4_(c0nm_headflit[4]), .c0nm_headflit_7_(c0nm_headflit[7]));
  /*CASIO@<instance>
     <id>mx387</id>
     <module>mux_merged_mx92</module>
     <compmap>F1:c0sm_b0m_v0m_u269, F2:c0sm_b0m_v0m_u268, F3:c0sm_b0m_v0m_u264, F4:c0sm_b0m_v0m_u263, F5:c0sm_b0m_v0m_u256, F6:c0sm_b0m_v0m_u255, F7:c0sm_b0m_v0m_u251, F8:c0sm_b0m_v0m_u250, F9:c0sm_b0m_v0m_u246, F10:c0sm_b0m_v0m_u245, F11:c0sm_b0m_v0m_u236, F12:c0sm_b0m_v0m_u235, F13:c0sm_b0m_v0m_u221, F14:c0sm_b0m_v0m_u220, F15:c0sm_b0m_v0m_u216, F16:c0sm_b0m_v0m_u215, F17:c0sm_b0m_v0m_u211, F18:c0sm_b0m_v0m_u210</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux_merged_mx92 mx387(.c0sm_b0m_v0m_buffers0_0_(c0sm_b0m_v0m_buffers0_0_), .c0sm_b0m_v0m_buffers0_10_(c0sm_b0m_v0m_buffers0_10_), .c0sm_b0m_v0m_buffers0_11_(c0sm_b0m_v0m_buffers0_11_), .c0sm_b0m_v0m_buffers0_1_(c0sm_b0m_v0m_buffers0_1_), .c0sm_b0m_v0m_buffers0_2_(c0sm_b0m_v0m_buffers0_2_), .c0sm_b0m_v0m_buffers0_4_(c0sm_b0m_v0m_buffers0_4_), .c0sm_b0m_v0m_buffers0_7_(c0sm_b0m_v0m_buffers0_7_), .c0sm_b0m_v0m_buffers0_8_(c0sm_b0m_v0m_buffers0_8_), .c0sm_b0m_v0m_buffers0_9_(c0sm_b0m_v0m_buffers0_9_), .c0sm_b0m_v0m_n105(c0sm_b0m_v0m_n105), .c0sm_b0m_v0m_n114(c0sm_b0m_v0m_n114), .c0sm_b0m_v0m_n122(c0sm_b0m_v0m_n122), .c0sm_b0m_v0m_n125(c0sm_b0m_v0m_n125), .c0sm_b0m_v0m_n131(c0sm_b0m_v0m_n131), .c0sm_b0m_v0m_n134(c0sm_b0m_v0m_n134), .c0sm_b0m_v0m_n144(c0sm_b0m_v0m_n144), .c0sm_b0m_v0m_n147(c0sm_b0m_v0m_n147), .c0sm_b0m_v0m_n162(c0sm_b0m_v0m_n162), .c0sm_b0m_v0m_n165(c0sm_b0m_v0m_n165), .c0sm_b0m_v0m_n168(c0sm_b0m_v0m_n168), .c0sm_b0m_v0m_n171(c0sm_b0m_v0m_n171), .c0sm_b0m_v0m_n174(c0sm_b0m_v0m_n174), .c0sm_b0m_v0m_n177(c0sm_b0m_v0m_n177), .c0sm_b0m_v0m_n180(c0sm_b0m_v0m_n180), .c0sm_b0m_v0m_n183(c0sm_b0m_v0m_n183), .c0sm_b0m_v0m_n186(c0sm_b0m_v0m_n186), .c0sm_b0m_v0m_n187(c0sm_b0m_v0m_n187), .c0sm_b0m_v0m_n190(c0sm_b0m_v0m_n190), .c0sm_b0m_v0m_n192(c0sm_b0m_v0m_n192), .c0sm_b0m_v0m_n193(c0sm_b0m_v0m_n193), .c0sm_b0m_v0m_n21(c0sm_b0m_v0m_n21), .c0sm_b0m_v0m_n23(c0sm_b0m_v0m_n23), .c0sm_b0m_v0m_n29(c0sm_b0m_v0m_n29), .c0sm_b0m_v0m_n35(c0sm_b0m_v0m_n35), .c0sm_b0m_v0m_n41(c0sm_b0m_v0m_n41), .c0sm_b0m_v0m_n62(c0sm_b0m_v0m_n62), .c0sm_b0m_v0m_n65(c0sm_b0m_v0m_n65), .c0sm_b0m_v0m_n68(c0sm_b0m_v0m_n68), .c0sm_b0m_v0m_n71(c0sm_b0m_v0m_n71), .c0sm_b0m_v0m_n73(c0sm_b0m_v0m_n73), .c0sm_b0m_headflit_10_(c0sm_b0m_headflit_10_), .c0sm_b0m_headflit_11_(c0sm_b0m_headflit_11_), .c0sm_b0m_headflit_8_(c0sm_b0m_headflit_8_), .c0sm_b0m_headflit_9_(c0sm_b0m_headflit_9_), .c0sm_headflit_0_(c0sm_headflit[0]), .c0sm_headflit_1_(c0sm_headflit[1]), .c0sm_headflit_2_(c0sm_headflit[2]), .c0sm_headflit_4_(c0sm_headflit[4]), .c0sm_headflit_7_(c0sm_headflit[7]));
  /*CASIO@<instance>
     <id>mx400</id>
     <module>mux_merged_mx93</module>
     <compmap>F1:c0nm_b0m_v0m_u268, F2:c0nm_b0m_v0m_u87, F3:c0nm_b0m_v0m_u86</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux_merged_mx93 mx400(.c0nm_b0m_v0m_buffers0_0_(c0nm_b0m_v0m_buffers0_0_), .c0nm_b0m_v0m_n105(c0nm_b0m_v0m_n105), .c0nm_b0m_v0m_n110(c0nm_b0m_v0m_n110), .c0nm_b0m_v0m_n111(c0nm_b0m_v0m_n111), .c0nm_b0m_v0m_n113(c0nm_b0m_v0m_n113), .c0nm_b0m_v0m_n114(c0nm_b0m_v0m_n114), .c0nm_b0m_v0m_n115(c0nm_b0m_v0m_n115), .c0nm_b0m_v0m_n187(c0nm_b0m_v0m_n187), .c0nm_b0m_v0m_n192(c0nm_b0m_v0m_n192), .c0nm_b0m_v0m_n193(c0nm_b0m_v0m_n193), .c0nm_b0m_v0m_n23(c0nm_b0m_v0m_n23), .c0nm_b0m_v0m_n276(c0nm_b0m_v0m_n276), .c0nm_b0m_v0m_n73(c0nm_b0m_v0m_n73), .debitout_0(debitout_0), .c0nm_b0m_v0m_n27(c0nm_b0m_v0m_n27), .c0nm_headflit_0_(c0nm_headflit[0]));
  /*CASIO@<instance>
     <id>mx401</id>
     <module>mux_merged_mx94</module>
     <compmap>F1:c0nm_b0m_v0m_u263, F2:c0nm_b0m_v0m_u94, F3:c0nm_b0m_v0m_u93</compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  mux_merged_mx94 mx401(.c0nm_b0m_v0m_buffers0_1_(c0nm_b0m_v0m_buffers0_1_), .c0nm_b0m_v0m_n110(c0nm_b0m_v0m_n110), .c0nm_b0m_v0m_n111(c0nm_b0m_v0m_n111), .c0nm_b0m_v0m_n113(c0nm_b0m_v0m_n113), .c0nm_b0m_v0m_n115(c0nm_b0m_v0m_n115), .c0nm_b0m_v0m_n122(c0nm_b0m_v0m_n122), .c0nm_b0m_v0m_n125(c0nm_b0m_v0m_n125), .c0nm_b0m_v0m_n187(c0nm_b0m_v0m_n187), .c0nm_b0m_v0m_n192(c0nm_b0m_v0m_n192), .c0nm_b0m_v0m_n193(c0nm_b0m_v0m_n193), .c0nm_b0m_v0m_n275(c0nm_b0m_v0m_n275), .c0nm_b0m_v0m_n29(c0nm_b0m_v0m_n29), .c0nm_b0m_v0m_n73(c0nm_b0m_v0m_n73), .debitout_0(debitout_0), .c0nm_b0m_v0m_n32(c0nm_b0m_v0m_n32), .c0nm_headflit_1_(c0nm_headflit[1]));
  /*CASIO@<instance>
     <id>mx404</id>
     <module>counter_mx95</module>
     <compmap>F1:c0nm_b0m_v0m_head_reg_1_, F2:c0nm_b0m_v0m_head_reg_0_, </compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  counter_mx95 mx404(.c0nm_b0m_v0m_n257(c0nm_b0m_v0m_n257), .c0nm_b0m_v0m_n258(c0nm_b0m_v0m_n258), .clk(clk), .c0nm_b0m_v0m_head_0_(c0nm_b0m_v0m_head_0_), .c0nm_b0m_v0m_head_1_(c0nm_b0m_v0m_head_1_));
  /*CASIO@<instance>
     <id>mx405</id>
     <module>counter_mx96</module>
     <compmap>F1:c0nm_b0m_v0m_tail_reg_0_, F2:c0nm_b0m_v0m_tail_reg_1_, </compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  counter_mx96 mx405(.c0nm_b0m_v0m_n260(c0nm_b0m_v0m_n260), .c0nm_b0m_v0m_n261(c0nm_b0m_v0m_n261), .clk(clk), .c0nm_b0m_v0m_tail_0_(c0nm_b0m_v0m_tail_0_), .c0nm_b0m_v0m_tail_1_(c0nm_b0m_v0m_tail_1_));
  /*CASIO@<instance>
     <id>mx406</id>
     <module>counter_mx97</module>
     <compmap>F1:c0sm_b0m_v0m_head_reg_1_, F2:c0sm_b0m_v0m_head_reg_0_, </compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  counter_mx97 mx406(.c0sm_b0m_v0m_n280(c0sm_b0m_v0m_n280), .c0sm_b0m_v0m_n281(c0sm_b0m_v0m_n281), .clk(clk), .c0sm_b0m_v0m_head_0_(c0sm_b0m_v0m_head_0_), .c0sm_b0m_v0m_head_1_(c0sm_b0m_v0m_head_1_));
  /*CASIO@<instance>
     <id>mx407</id>
     <module>counter_mx98</module>
     <compmap>F1:c0sm_b0m_v0m_tail_reg_0_, F2:c0sm_b0m_v0m_tail_reg_1_, </compmap>
     <creationtool>bsim</creationtool>
     <confidence>0.60</confidence>
     <flag></flag>
     <wiremap></wiremap>
     </instance>
   */
  counter_mx98 mx407(.c0sm_b0m_v0m_n277(c0sm_b0m_v0m_n277), .c0sm_b0m_v0m_n278(c0sm_b0m_v0m_n278), .clk(clk), .c0sm_b0m_v0m_tail_0_(c0sm_b0m_v0m_tail_0_), .c0sm_b0m_v0m_tail_1_(c0sm_b0m_v0m_tail_1_));
endmodule
