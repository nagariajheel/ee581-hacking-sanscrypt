module mux21_mx0 
(
  s0m_m0m_n1, 
  s0m_m0m_row1_0_, 
  s0m_request1_0_, 
  s0m_m0m_n2,
  s0m_m0m_n3
);
  input s0m_m0m_n1;
  input s0m_m0m_row1_0_;
  input s0m_request1_0_;
  output s0m_m0m_n2;
  output s0m_m0m_n3;
  wire s0m__logic0_;
  wire s0m_outb0_0_;

  // moduleNum: x0
  // type: mux21
  // conflicting modules: 
  // number of bit inputs: 1
  // number of bit outputs: 0
  // number of word inputs: 2
  // number of word outputs: 1
  // number of internal gates: 4
  // number of non-inferred gates: 0
  // ILP vars: 21/23
  // type: INFERRED
  // marked bad? no
  // input word of size 2 : index:6 s0m_m0m_n1 s0m_m0m_n1 
  // input word of size 2 : index:7 s0m_request1[0] s0m_request1[0] 
  // output word of size 2 : index:8 s0m_m0m_n3 s0m_m0m_n2 
  // group: sel; nodes: [ s0m_m0m_row1_0_ ]

  TIELO_X1M_A12TR s0m_u2 (.Y(s0m__logic0_));
  AOI21_X0P5M_A12TR s0m_m0m_u7 (.A0(s0m_request1_0_), .A1(s0m_m0m_row1_0_), .B0(s0m_m0m_n1), .Y(s0m_outb0_0_));
  AOI2XB1_X0P5M_A12TR s0m_m0m_u6 (.A0(s0m_m0m_row1_0_), .A1N(s0m_request1_0_), .B0(s0m_outb0_0_), .Y(s0m_m0m_n3));
  XOR2_X0P5M_A12TR s0m_m0m_u5 (.A(s0m__logic0_), .B(s0m_m0m_n3), .Y(s0m_m0m_n2));
endmodule
module mux21_mx1 
(
  flitout_switch_0_0_, 
  flitout_switch_0_11_, 
  flitout_switch_0_1_, 
  flitout_switch_0_4_, 
  flitout_switch_1_0_, 
  flitout_switch_1_11_, 
  flitout_switch_1_1_, 
  flitout_switch_1_4_, 
  x0m_colsel1reg_0_, 
  x0m_bx0m_m1m_int01,
  x0m_bx11m_m1m_int01,
  x0m_bx1m_m1m_int01,
  x0m_bx4m_m1m_int01
);
  input flitout_switch_0_0_;
  input flitout_switch_0_11_;
  input flitout_switch_0_1_;
  input flitout_switch_0_4_;
  input flitout_switch_1_0_;
  input flitout_switch_1_11_;
  input flitout_switch_1_1_;
  input flitout_switch_1_4_;
  input x0m_colsel1reg_0_;
  output x0m_bx0m_m1m_int01;
  output x0m_bx11m_m1m_int01;
  output x0m_bx1m_m1m_int01;
  output x0m_bx4m_m1m_int01;

  // moduleNum: x1
  // type: mux21
  // conflicting modules: 
  // number of bit inputs: 1
  // number of bit outputs: 0
  // number of word inputs: 2
  // number of word outputs: 1
  // number of internal gates: 4
  // number of non-inferred gates: 0
  // ILP vars: 53/64
  // type: INFERRED
  // marked bad? no
  // input word of size 4 : index:-1 flitout_switch_0[4] flitout_switch_0[0] flitout_switch_0[11] flitout_switch_0[1] 
  // input word of size 4 : index:-1 flitout_switch_1[4] flitout_switch_1[0] flitout_switch_1[11] flitout_switch_1[1] 
  // output word of size 4 : index:238 x0m_bx4m_m1m_int01 x0m_bx0m_m1m_int01 x0m_bx11m_m1m_int01 x0m_bx1m_m1m_int01 
  // group: sel; nodes: [ x0m_colsel1reg_0_ ]

  MXT2_X0P5M_A12TR x0m_bx0m_m1m_m0m_u1 (.A(flitout_switch_0_0_), .B(flitout_switch_1_0_), .S0(x0m_colsel1reg_0_), .Y(x0m_bx0m_m1m_int01));
  MXT2_X0P5M_A12TR x0m_bx1m_m1m_m0m_u1 (.A(flitout_switch_0_1_), .B(flitout_switch_1_1_), .S0(x0m_colsel1reg_0_), .Y(x0m_bx1m_m1m_int01));
  MXT2_X0P5M_A12TR x0m_bx4m_m1m_m0m_u1 (.A(flitout_switch_0_4_), .B(flitout_switch_1_4_), .S0(x0m_colsel1reg_0_), .Y(x0m_bx4m_m1m_int01));
  MXT2_X0P5M_A12TR x0m_bx11m_m1m_m0m_u1 (.A(flitout_switch_0_11_), .B(flitout_switch_1_11_), .S0(x0m_colsel1reg_0_), .Y(x0m_bx11m_m1m_int01));
endmodule
module mux21_mx2 
(
  x0m__logic0_, 
  x0m_bx11m_m1m_int01, 
  x0m_bx4m_m1m_int01, 
  x0m_colsel1reg_1_, 
  flitout_1_11_,
  flitout_1_4_
);
  input x0m__logic0_;
  input x0m_bx11m_m1m_int01;
  input x0m_bx4m_m1m_int01;
  input x0m_colsel1reg_1_;
  output flitout_1_11_;
  output flitout_1_4_;

  // moduleNum: x2
  // type: mux21
  // conflicting modules: 
  // number of bit inputs: 1
  // number of bit outputs: 0
  // number of word inputs: 2
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 65/77
  // type: INFERRED
  // marked bad? no
  // input word of size 2 : index:-1 x0m_bx11m_m1m_int01 x0m_bx4m_m1m_int01 
  // input word of size 10 : index:-1 x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_
  // x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_
  // output word of size 2 : index:239 flitout_1[11] flitout_1[4] 
  // group: sel; nodes: [ x0m_colsel1reg_1_ ]

  MXT2_X0P5M_A12TR x0m_bx4m_m1m_m4m_u1 (.A(x0m_bx4m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1_4_));
  MXT2_X0P5M_A12TR x0m_bx11m_m1m_m4m_u1 (.A(x0m_bx11m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1_11_));
endmodule
module mux21i_mx3 
(
  c0nm_routewire_0_, 
  c0nm_routewire_1_, 
  c0nm_v0m_n3, 
  c0nm_v0m_n4, 
  c0nm_v0m_n7, 
  c0nm_v0m_n2,
  c0nm_v0m_n6
);
  input c0nm_routewire_0_;
  input c0nm_routewire_1_;
  input c0nm_v0m_n3;
  input c0nm_v0m_n4;
  input c0nm_v0m_n7;
  output c0nm_v0m_n2;
  output c0nm_v0m_n6;

  // moduleNum: x3
  // type: mux21i
  // conflicting modules: 
  // number of bit inputs: 1
  // number of bit outputs: 0
  // number of word inputs: 2
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 90/90
  // type: INFERRED
  // marked bad? no
  // input word of size 2 : index:36 c0nm_v0m_n7 c0nm_v0m_n3 
  // input word of size 2 : index:37 c0nm_routewire[0] c0nm_routewire[1] 
  // output word of size 2 : index:38 c0nm_v0m_n6 c0nm_v0m_n2 
  // group: sel; nodes: [ c0nm_v0m_n4 ]

  MXIT2_X0P5M_A12TR c0nm_v0m_u7 (.A(c0nm_v0m_n7), .B(c0nm_routewire_0_), .S0(c0nm_v0m_n4), .Y(c0nm_v0m_n6));
  MXIT2_X0P5M_A12TR c0nm_v0m_u4 (.A(c0nm_v0m_n3), .B(c0nm_routewire_1_), .S0(c0nm_v0m_n4), .Y(c0nm_v0m_n2));
endmodule
module mux21i_mx4 
(
  c0nm_v0m_n18, 
  c0nm_v0m_n20, 
  c0nm_v0m_n21, 
  c0nm_v0m_state_queuelen_0_, 
  c0nm_v0m_state_queuelen_1_, 
  c0nm_v0m_n15,
  c0nm_v0m_n19
);
  input c0nm_v0m_n18;
  input c0nm_v0m_n20;
  input c0nm_v0m_n21;
  input c0nm_v0m_state_queuelen_0_;
  input c0nm_v0m_state_queuelen_1_;
  output c0nm_v0m_n15;
  output c0nm_v0m_n19;

  // moduleNum: x4
  // type: mux21i
  // conflicting modules: 
  // number of bit inputs: 1
  // number of bit outputs: 0
  // number of word inputs: 2
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 91/91
  // type: INFERRED
  // marked bad? no
  // input word of size 2 : index:39 c0nm_v0m_state_queuelen_0_ c0nm_v0m_n20 
  // input word of size 2 : index:40 c0nm_v0m_n18 c0nm_v0m_n21 
  // output word of size 2 : index:41 c0nm_v0m_n15 c0nm_v0m_n19 
  // group: sel; nodes: [ c0nm_v0m_state_queuelen_1_ ]

  MXIT2_X0P5M_A12TR c0nm_v0m_u18 (.A(c0nm_v0m_n20), .B(c0nm_v0m_n21), .S0(c0nm_v0m_state_queuelen_1_), .Y(c0nm_v0m_n19));
  MXIT2_X0P5M_A12TR c0nm_v0m_u16 (.A(c0nm_v0m_state_queuelen_0_), .B(c0nm_v0m_n18), .S0(c0nm_v0m_state_queuelen_1_), .Y(c0nm_v0m_n15));
endmodule
module mux21i_mx5 
(
  c0sm_routewire_0_, 
  c0sm_routewire_1_, 
  c0sm_v0m_n3, 
  c0sm_v0m_n4, 
  c0sm_v0m_n7, 
  c0sm_v0m_n2,
  c0sm_v0m_n6
);
  input c0sm_routewire_0_;
  input c0sm_routewire_1_;
  input c0sm_v0m_n3;
  input c0sm_v0m_n4;
  input c0sm_v0m_n7;
  output c0sm_v0m_n2;
  output c0sm_v0m_n6;

  // moduleNum: x5
  // type: mux21i
  // conflicting modules: 
  // number of bit inputs: 1
  // number of bit outputs: 0
  // number of word inputs: 2
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 104/104
  // type: INFERRED
  // marked bad? no
  // input word of size 2 : index:54 c0sm_v0m_n7 c0sm_v0m_n3 
  // input word of size 2 : index:55 c0sm_routewire[0] c0sm_routewire[1] 
  // output word of size 2 : index:56 c0sm_v0m_n6 c0sm_v0m_n2 
  // group: sel; nodes: [ c0sm_v0m_n4 ]

  MXIT2_X0P5M_A12TR c0sm_v0m_u7 (.A(c0sm_v0m_n7), .B(c0sm_routewire_0_), .S0(c0sm_v0m_n4), .Y(c0sm_v0m_n6));
  MXIT2_X0P5M_A12TR c0sm_v0m_u4 (.A(c0sm_v0m_n3), .B(c0sm_routewire_1_), .S0(c0sm_v0m_n4), .Y(c0sm_v0m_n2));
endmodule
module mux21i_mx6 
(
  c0sm_v0m_n18, 
  c0sm_v0m_n20, 
  c0sm_v0m_n21, 
  c0sm_v0m_state_queuelen_0_, 
  c0sm_v0m_state_queuelen_1_, 
  c0sm_v0m_n15,
  c0sm_v0m_n19
);
  input c0sm_v0m_n18;
  input c0sm_v0m_n20;
  input c0sm_v0m_n21;
  input c0sm_v0m_state_queuelen_0_;
  input c0sm_v0m_state_queuelen_1_;
  output c0sm_v0m_n15;
  output c0sm_v0m_n19;

  // moduleNum: x6
  // type: mux21i
  // conflicting modules: 
  // number of bit inputs: 1
  // number of bit outputs: 0
  // number of word inputs: 2
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 105/105
  // type: INFERRED
  // marked bad? no
  // input word of size 2 : index:57 c0sm_v0m_state_queuelen_0_ c0sm_v0m_n20 
  // input word of size 2 : index:58 c0sm_v0m_n18 c0sm_v0m_n21 
  // output word of size 2 : index:59 c0sm_v0m_n15 c0sm_v0m_n19 
  // group: sel; nodes: [ c0sm_v0m_state_queuelen_1_ ]

  MXIT2_X0P5M_A12TR c0sm_v0m_u18 (.A(c0sm_v0m_n20), .B(c0sm_v0m_n21), .S0(c0sm_v0m_state_queuelen_1_), .Y(c0sm_v0m_n19));
  MXIT2_X0P5M_A12TR c0sm_v0m_u16 (.A(c0sm_v0m_state_queuelen_0_), .B(c0sm_v0m_n18), .S0(c0sm_v0m_state_queuelen_1_), .Y(c0sm_v0m_n15));
endmodule
module mux21i_mx7 
(
  s0m_n13, 
  s0m_n14, 
  s0m_n15, 
  s0m_n17, 
  s0m_n18, 
  s0m_n22,
  s0m_n23
);
  input s0m_n13;
  input s0m_n14;
  input s0m_n15;
  input s0m_n17;
  input s0m_n18;
  output s0m_n22;
  output s0m_n23;

  // moduleNum: x7
  // type: mux21i
  // conflicting modules: 
  // number of bit inputs: 1
  // number of bit outputs: 0
  // number of word inputs: 2
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 106/106
  // type: INFERRED
  // marked bad? no
  // input word of size 2 : index:60 s0m_n13 s0m_n17 
  // input word of size 2 : index:61 s0m_n14 s0m_n18 
  // output word of size 2 : index:62 s0m_n23 s0m_n22 
  // group: sel; nodes: [ s0m_n15 ]

  MXIT2_X0P5M_A12TR s0m_u28 (.A(s0m_n17), .B(s0m_n18), .S0(s0m_n15), .Y(s0m_n22));
  MXIT2_X0P5M_A12TR s0m_u25 (.A(s0m_n13), .B(s0m_n14), .S0(s0m_n15), .Y(s0m_n23));
endmodule
module mux21i_mx8 
(
  s0m_n10, 
  s0m_n11, 
  s0m_n6, 
  s0m_n7, 
  s0m_n8, 
  s0m_n24,
  s0m_n25
);
  input s0m_n10;
  input s0m_n11;
  input s0m_n6;
  input s0m_n7;
  input s0m_n8;
  output s0m_n24;
  output s0m_n25;

  // moduleNum: x8
  // type: mux21i
  // conflicting modules: 
  // number of bit inputs: 1
  // number of bit outputs: 0
  // number of word inputs: 2
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 107/107
  // type: INFERRED
  // marked bad? no
  // input word of size 2 : index:63 s0m_n6 s0m_n10 
  // input word of size 2 : index:64 s0m_n7 s0m_n11 
  // output word of size 2 : index:65 s0m_n25 s0m_n24 
  // group: sel; nodes: [ s0m_n8 ]

  MXIT2_X0P5M_A12TR s0m_u19 (.A(s0m_n10), .B(s0m_n11), .S0(s0m_n8), .Y(s0m_n24));
  MXIT2_X0P5M_A12TR s0m_u16 (.A(s0m_n6), .B(s0m_n7), .S0(s0m_n8), .Y(s0m_n25));
endmodule
module mux21i_mx9 
(
  c0nm_v0m_n9, 
  s0m_n26, 
  s0m_n4, 
  s0m_n5, 
  s0m_state_invc0_0_, 
  nomorebufs_0,
  s0m_debit_outvc0
);
  input c0nm_v0m_n9;
  input s0m_n26;
  input s0m_n4;
  input s0m_n5;
  input s0m_state_invc0_0_;
  output nomorebufs_0;
  output s0m_debit_outvc0;

  // moduleNum: x9
  // type: mux21i
  // conflicting modules: 
  // number of bit inputs: 1
  // number of bit outputs: 0
  // number of word inputs: 2
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 108/108
  // type: INFERRED
  // marked bad? no
  // input word of size 2 : index:66 s0m_n4 s0m_n26 
  // input word of size 2 : index:67 s0m_n5 c0nm_v0m_n9 
  // output word of size 2 : index:68 nomorebufs_0 s0m_debit_outvc0 
  // group: sel; nodes: [ s0m_state_invc0_0_ ]

  MXIT2_X0P5M_A12TR s0m_u36 (.A(s0m_n26), .B(c0nm_v0m_n9), .S0(s0m_state_invc0_0_), .Y(s0m_debit_outvc0));
  MXIT2_X0P5M_A12TR s0m_u13 (.A(s0m_n4), .B(s0m_n5), .S0(s0m_state_invc0_0_), .Y(nomorebufs_0));
endmodule
module mux21i_mx10 
(
  c0nm_v0m_n9, 
  s0m_n1, 
  s0m_n2, 
  s0m_n20, 
  s0m_state_invc1_0_, 
  s0m_debit_outvc1,
  s0m_tail_outvc1
);
  input c0nm_v0m_n9;
  input s0m_n1;
  input s0m_n2;
  input s0m_n20;
  input s0m_state_invc1_0_;
  output s0m_debit_outvc1;
  output s0m_tail_outvc1;

  // moduleNum: x10
  // type: mux21i
  // conflicting modules: 
  // number of bit inputs: 1
  // number of bit outputs: 0
  // number of word inputs: 2
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 109/109
  // type: INFERRED
  // marked bad? no
  // input word of size 2 : index:69 s0m_n1 s0m_n20 
  // input word of size 2 : index:70 s0m_n2 c0nm_v0m_n9 
  // output word of size 2 : index:71 s0m_tail_outvc1 s0m_debit_outvc1 
  // group: sel; nodes: [ s0m_state_invc1_0_ ]

  MXIT2_X0P5M_A12TR s0m_u34 (.A(s0m_n20), .B(c0nm_v0m_n9), .S0(s0m_state_invc1_0_), .Y(s0m_debit_outvc1));
  MXIT2_X0P5M_A12TR s0m_u3 (.A(s0m_n1), .B(s0m_n2), .S0(s0m_state_invc1_0_), .Y(s0m_tail_outvc1));
endmodule
module mux21i_aoi22_mx11 
(
  c0nm_r0m_n13, 
  c0nm_r0m_n14, 
  c0sm_r0m_n13, 
  c0sm_r0m_n14, 
  curry_0_, 
  curry_1_, 
  c0nm_r0m_n12,
  c0sm_r0m_n12
);
  input c0nm_r0m_n13;
  input c0nm_r0m_n14;
  input c0sm_r0m_n13;
  input c0sm_r0m_n14;
  input curry_0_;
  input curry_1_;
  output c0nm_r0m_n12;
  output c0sm_r0m_n12;

  // moduleNum: x11
  // type: mux21i_aoi22
  // conflicting modules: 
  // number of bit inputs: 6
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 132/132
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:74 c0nm_r0m_n12 c0sm_r0m_n12 
  // group: sel; nodes: [ curry[1] curry[0] ]

  AOI22_X0P5M_A12TR c0nm_r0m_u12 (.A0(c0nm_r0m_n13), .A1(curry_0_), .B0(curry_1_), .B1(c0nm_r0m_n14), .Y(c0nm_r0m_n12));
  AOI22_X0P5M_A12TR c0sm_r0m_u12 (.A0(c0sm_r0m_n13), .A1(curry_0_), .B0(curry_1_), .B1(c0sm_r0m_n14), .Y(c0sm_r0m_n12));
endmodule
module mux21i_aoi22_mx12 
(
  c0nm_b0m_n1, 
  c0nm_b0m_v0m_n114, 
  c0nm_b0m_v0m_n119, 
  c0nm_b0m_v0m_n125, 
  flitin_0_0_, 
  flitin_0_1_, 
  c0nm_b0m_v0m_n118,
  c0nm_b0m_v0m_n127
);
  input c0nm_b0m_n1;
  input c0nm_b0m_v0m_n114;
  input c0nm_b0m_v0m_n119;
  input c0nm_b0m_v0m_n125;
  input flitin_0_0_;
  input flitin_0_1_;
  output c0nm_b0m_v0m_n118;
  output c0nm_b0m_v0m_n127;

  // moduleNum: x12
  // type: mux21i_aoi22
  // conflicting modules: 
  // number of bit inputs: 6
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 133/133
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:75 c0nm_b0m_v0m_n127 c0nm_b0m_v0m_n118 
  // group: sel; nodes: [ c0nm_b0m_n1 c0nm_b0m_v0m_n119 ]

  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u96 (.A0(c0nm_b0m_v0m_n119), .A1(c0nm_b0m_v0m_n125), .B0(flitin_0_1_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n127));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u89 (.A0(c0nm_b0m_v0m_n119), .A1(c0nm_b0m_v0m_n114), .B0(flitin_0_0_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n118));
endmodule
module mux21i_aoi22_mx13 
(
  c0nm_b0m_n1, 
  c0nm_b0m_v0m_buffers3_10_, 
  c0nm_b0m_v0m_buffers3_11_, 
  c0nm_b0m_v0m_buffers3_2_, 
  c0nm_b0m_v0m_buffers3_3_, 
  c0nm_b0m_v0m_buffers3_4_, 
  c0nm_b0m_v0m_buffers3_5_, 
  c0nm_b0m_v0m_buffers3_6_, 
  c0nm_b0m_v0m_buffers3_7_, 
  c0nm_b0m_v0m_buffers3_8_, 
  c0nm_b0m_v0m_buffers3_9_, 
  c0nm_b0m_v0m_n128, 
  c0nm_b0m_wdata_10_, 
  c0nm_b0m_wdata_11_, 
  c0nm_b0m_wdata_2_, 
  c0nm_b0m_wdata_3_, 
  c0nm_b0m_wdata_4_, 
  c0nm_b0m_wdata_5_, 
  c0nm_b0m_wdata_6_, 
  c0nm_b0m_wdata_7_, 
  c0nm_b0m_wdata_8_, 
  c0nm_b0m_wdata_9_, 
  flitin_0_10_, 
  flitin_0_11_, 
  flitin_0_2_, 
  flitin_0_3_, 
  flitin_0_4_, 
  flitin_0_5_, 
  flitin_0_6_, 
  flitin_0_7_, 
  flitin_0_8_, 
  flitin_0_9_, 
  c0nm_b0m_v0m_n137,
  c0nm_b0m_v0m_n143,
  c0nm_b0m_v0m_n149,
  c0nm_b0m_v0m_n155,
  c0nm_b0m_v0m_n161,
  c0nm_b0m_v0m_n167,
  c0nm_b0m_v0m_n173,
  c0nm_b0m_v0m_n179,
  c0nm_b0m_v0m_n185,
  c0nm_b0m_v0m_n195
);
  input c0nm_b0m_n1;
  input c0nm_b0m_v0m_buffers3_10_;
  input c0nm_b0m_v0m_buffers3_11_;
  input c0nm_b0m_v0m_buffers3_2_;
  input c0nm_b0m_v0m_buffers3_3_;
  input c0nm_b0m_v0m_buffers3_4_;
  input c0nm_b0m_v0m_buffers3_5_;
  input c0nm_b0m_v0m_buffers3_6_;
  input c0nm_b0m_v0m_buffers3_7_;
  input c0nm_b0m_v0m_buffers3_8_;
  input c0nm_b0m_v0m_buffers3_9_;
  input c0nm_b0m_v0m_n128;
  input c0nm_b0m_wdata_10_;
  input c0nm_b0m_wdata_11_;
  input c0nm_b0m_wdata_2_;
  input c0nm_b0m_wdata_3_;
  input c0nm_b0m_wdata_4_;
  input c0nm_b0m_wdata_5_;
  input c0nm_b0m_wdata_6_;
  input c0nm_b0m_wdata_7_;
  input c0nm_b0m_wdata_8_;
  input c0nm_b0m_wdata_9_;
  input flitin_0_10_;
  input flitin_0_11_;
  input flitin_0_2_;
  input flitin_0_3_;
  input flitin_0_4_;
  input flitin_0_5_;
  input flitin_0_6_;
  input flitin_0_7_;
  input flitin_0_8_;
  input flitin_0_9_;
  output c0nm_b0m_v0m_n137;
  output c0nm_b0m_v0m_n143;
  output c0nm_b0m_v0m_n149;
  output c0nm_b0m_v0m_n155;
  output c0nm_b0m_v0m_n161;
  output c0nm_b0m_v0m_n167;
  output c0nm_b0m_v0m_n173;
  output c0nm_b0m_v0m_n179;
  output c0nm_b0m_v0m_n185;
  output c0nm_b0m_v0m_n195;

  // moduleNum: x13
  // type: mux21i_aoi22
  // conflicting modules: 
  // number of bit inputs: 32
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 134/154
  // type: INFERRED
  // marked bad? no
  // output word of size 20 : index:76 c0nm_b0m_v0m_n137 c0nm_b0m_v0m_n137 c0nm_b0m_v0m_n143 c0nm_b0m_v0m_n143
  // c0nm_b0m_v0m_n185 c0nm_b0m_v0m_n185 c0nm_b0m_v0m_n167 c0nm_b0m_v0m_n167 c0nm_b0m_v0m_n173 c0nm_b0m_v0m_n173
  // c0nm_b0m_v0m_n179 c0nm_b0m_v0m_n179 c0nm_b0m_v0m_n161 c0nm_b0m_v0m_n161 c0nm_b0m_v0m_n155 c0nm_b0m_v0m_n155
  // c0nm_b0m_v0m_n149 c0nm_b0m_v0m_n149 c0nm_b0m_v0m_n195 c0nm_b0m_v0m_n195
  // group: sel; nodes: [ c0nm_b0m_n1 c0nm_b0m_v0m_n128 ]

  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u181 (.A0(c0nm_b0m_v0m_buffers3_11_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_n1), .B1(c0nm_b0m_wdata_11_), .Y(c0nm_b0m_v0m_n195));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u160 (.A0(c0nm_b0m_v0m_buffers3_10_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_10_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n185));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u153 (.A0(c0nm_b0m_v0m_buffers3_9_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_9_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n179));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u146 (.A0(c0nm_b0m_v0m_buffers3_8_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_8_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n173));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u139 (.A0(c0nm_b0m_v0m_buffers3_7_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_7_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n167));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u132 (.A0(c0nm_b0m_v0m_buffers3_6_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_6_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n161));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u125 (.A0(c0nm_b0m_v0m_buffers3_5_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_5_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n155));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u118 (.A0(c0nm_b0m_v0m_buffers3_4_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_4_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n149));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u111 (.A0(c0nm_b0m_v0m_buffers3_3_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_3_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n143));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u104 (.A0(c0nm_b0m_v0m_buffers3_2_), .A1(c0nm_b0m_v0m_n128), .B0(c0nm_b0m_wdata_2_), .B1(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n137));
endmodule
module mux21i_aoi22_mx14 
(
  c0nm_b0m_v0m_buffers0_0_, 
  c0nm_b0m_v0m_buffers0_1_, 
  c0nm_b0m_v0m_buffers0_3_, 
  c0nm_b0m_v0m_buffers0_5_, 
  c0nm_b0m_v0m_buffers0_6_, 
  c0nm_b0m_v0m_n114, 
  c0nm_b0m_v0m_n125, 
  c0nm_b0m_v0m_n141, 
  c0nm_b0m_v0m_n153, 
  c0nm_b0m_v0m_n159, 
  c0nm_b0m_v0m_n192, 
  c0nm_b0m_v0m_n193, 
  c0nm_b0m_v0m_n268,
  c0nm_b0m_v0m_n269,
  c0nm_b0m_v0m_n271,
  c0nm_b0m_v0m_n275,
  c0nm_b0m_v0m_n276
);
  input c0nm_b0m_v0m_buffers0_0_;
  input c0nm_b0m_v0m_buffers0_1_;
  input c0nm_b0m_v0m_buffers0_3_;
  input c0nm_b0m_v0m_buffers0_5_;
  input c0nm_b0m_v0m_buffers0_6_;
  input c0nm_b0m_v0m_n114;
  input c0nm_b0m_v0m_n125;
  input c0nm_b0m_v0m_n141;
  input c0nm_b0m_v0m_n153;
  input c0nm_b0m_v0m_n159;
  input c0nm_b0m_v0m_n192;
  input c0nm_b0m_v0m_n193;
  output c0nm_b0m_v0m_n268;
  output c0nm_b0m_v0m_n269;
  output c0nm_b0m_v0m_n271;
  output c0nm_b0m_v0m_n275;
  output c0nm_b0m_v0m_n276;

  // moduleNum: x14
  // type: mux21i_aoi22
  // conflicting modules: 
  // number of bit inputs: 12
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 5
  // number of non-inferred gates: 0
  // ILP vars: 185/197
  // type: INFERRED
  // marked bad? no
  // output word of size 5 : index:240 c0nm_b0m_v0m_n269 c0nm_b0m_v0m_n268 c0nm_b0m_v0m_n276 c0nm_b0m_v0m_n275
  // c0nm_b0m_v0m_n271
  // group: sel; nodes: [ c0nm_b0m_v0m_n193 c0nm_b0m_v0m_n192 ]

  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u269 (.A0(c0nm_b0m_v0m_buffers0_0_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n114), .Y(c0nm_b0m_v0m_n276));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u264 (.A0(c0nm_b0m_v0m_buffers0_1_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n125), .Y(c0nm_b0m_v0m_n275));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u241 (.A0(c0nm_b0m_v0m_buffers0_3_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n141), .Y(c0nm_b0m_v0m_n271));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u231 (.A0(c0nm_b0m_v0m_buffers0_5_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n153), .Y(c0nm_b0m_v0m_n269));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u226 (.A0(c0nm_b0m_v0m_buffers0_6_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n159), .Y(c0nm_b0m_v0m_n268));
endmodule
module mux21i_aoi22_mx15 
(
  c0nm_b0m_v0m_buffers0_0_, 
  c0nm_b0m_v0m_buffers0_10_, 
  c0nm_b0m_v0m_buffers0_11_, 
  c0nm_b0m_v0m_buffers0_1_, 
  c0nm_b0m_v0m_buffers0_2_, 
  c0nm_b0m_v0m_buffers0_3_, 
  c0nm_b0m_v0m_buffers0_4_, 
  c0nm_b0m_v0m_buffers0_5_, 
  c0nm_b0m_v0m_buffers0_6_, 
  c0nm_b0m_v0m_buffers0_7_, 
  c0nm_b0m_v0m_buffers0_8_, 
  c0nm_b0m_v0m_buffers0_9_, 
  c0nm_b0m_v0m_buffers2_0_, 
  c0nm_b0m_v0m_buffers2_10_, 
  c0nm_b0m_v0m_buffers2_11_, 
  c0nm_b0m_v0m_buffers2_1_, 
  c0nm_b0m_v0m_buffers2_2_, 
  c0nm_b0m_v0m_buffers2_3_, 
  c0nm_b0m_v0m_buffers2_4_, 
  c0nm_b0m_v0m_buffers2_5_, 
  c0nm_b0m_v0m_buffers2_6_, 
  c0nm_b0m_v0m_buffers2_7_, 
  c0nm_b0m_v0m_buffers2_8_, 
  c0nm_b0m_v0m_buffers2_9_, 
  c0nm_b0m_v0m_n120, 
  c0nm_b0m_v0m_n121, 
  c0nm_b0m_v0m_n117,
  c0nm_b0m_v0m_n126,
  c0nm_b0m_v0m_n136,
  c0nm_b0m_v0m_n142,
  c0nm_b0m_v0m_n148,
  c0nm_b0m_v0m_n154,
  c0nm_b0m_v0m_n160,
  c0nm_b0m_v0m_n166,
  c0nm_b0m_v0m_n172,
  c0nm_b0m_v0m_n178,
  c0nm_b0m_v0m_n184,
  c0nm_b0m_v0m_n194
);
  input c0nm_b0m_v0m_buffers0_0_;
  input c0nm_b0m_v0m_buffers0_10_;
  input c0nm_b0m_v0m_buffers0_11_;
  input c0nm_b0m_v0m_buffers0_1_;
  input c0nm_b0m_v0m_buffers0_2_;
  input c0nm_b0m_v0m_buffers0_3_;
  input c0nm_b0m_v0m_buffers0_4_;
  input c0nm_b0m_v0m_buffers0_5_;
  input c0nm_b0m_v0m_buffers0_6_;
  input c0nm_b0m_v0m_buffers0_7_;
  input c0nm_b0m_v0m_buffers0_8_;
  input c0nm_b0m_v0m_buffers0_9_;
  input c0nm_b0m_v0m_buffers2_0_;
  input c0nm_b0m_v0m_buffers2_10_;
  input c0nm_b0m_v0m_buffers2_11_;
  input c0nm_b0m_v0m_buffers2_1_;
  input c0nm_b0m_v0m_buffers2_2_;
  input c0nm_b0m_v0m_buffers2_3_;
  input c0nm_b0m_v0m_buffers2_4_;
  input c0nm_b0m_v0m_buffers2_5_;
  input c0nm_b0m_v0m_buffers2_6_;
  input c0nm_b0m_v0m_buffers2_7_;
  input c0nm_b0m_v0m_buffers2_8_;
  input c0nm_b0m_v0m_buffers2_9_;
  input c0nm_b0m_v0m_n120;
  input c0nm_b0m_v0m_n121;
  output c0nm_b0m_v0m_n117;
  output c0nm_b0m_v0m_n126;
  output c0nm_b0m_v0m_n136;
  output c0nm_b0m_v0m_n142;
  output c0nm_b0m_v0m_n148;
  output c0nm_b0m_v0m_n154;
  output c0nm_b0m_v0m_n160;
  output c0nm_b0m_v0m_n166;
  output c0nm_b0m_v0m_n172;
  output c0nm_b0m_v0m_n178;
  output c0nm_b0m_v0m_n184;
  output c0nm_b0m_v0m_n194;

  // moduleNum: x15
  // type: mux21i_aoi22
  // conflicting modules: 
  // number of bit inputs: 26
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 12
  // number of non-inferred gates: 0
  // ILP vars: 228/240
  // type: INFERRED
  // marked bad? no
  // output word of size 12 : index:98 c0nm_b0m_v0m_n172 c0nm_b0m_v0m_n126 c0nm_b0m_v0m_n178 c0nm_b0m_v0m_n184
  // c0nm_b0m_v0m_n117 c0nm_b0m_v0m_n194 c0nm_b0m_v0m_n154 c0nm_b0m_v0m_n160 c0nm_b0m_v0m_n142 c0nm_b0m_v0m_n166
  // c0nm_b0m_v0m_n136 c0nm_b0m_v0m_n148
  // group: sel; nodes: [ c0nm_b0m_v0m_n121 c0nm_b0m_v0m_n120 ]

  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u184 (.A0(c0nm_b0m_v0m_buffers2_11_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_11_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n194));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u161 (.A0(c0nm_b0m_v0m_buffers2_10_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_10_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n184));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u154 (.A0(c0nm_b0m_v0m_buffers2_9_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_9_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n178));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u147 (.A0(c0nm_b0m_v0m_buffers2_8_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_8_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n172));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u140 (.A0(c0nm_b0m_v0m_buffers2_7_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_7_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n166));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u133 (.A0(c0nm_b0m_v0m_buffers2_6_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_6_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n160));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u126 (.A0(c0nm_b0m_v0m_buffers2_5_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_5_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n154));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u119 (.A0(c0nm_b0m_v0m_buffers2_4_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_4_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n148));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u112 (.A0(c0nm_b0m_v0m_buffers2_3_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_3_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n142));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u105 (.A0(c0nm_b0m_v0m_buffers2_2_), .A1(c0nm_b0m_v0m_n121), .B0(c0nm_b0m_v0m_buffers0_2_), .B1(c0nm_b0m_v0m_n120), .Y(c0nm_b0m_v0m_n136));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u97 (.A0(c0nm_b0m_v0m_buffers0_1_), .A1(c0nm_b0m_v0m_n120), .B0(c0nm_b0m_v0m_buffers2_1_), .B1(c0nm_b0m_v0m_n121), .Y(c0nm_b0m_v0m_n126));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u90 (.A0(c0nm_b0m_v0m_buffers0_0_), .A1(c0nm_b0m_v0m_n120), .B0(c0nm_b0m_v0m_buffers2_0_), .B1(c0nm_b0m_v0m_n121), .Y(c0nm_b0m_v0m_n117));
endmodule
module mux21i_aoi22_mx16 
(
  c0nm_b0m_v0m_buffers0_10_, 
  c0nm_b0m_v0m_buffers0_11_, 
  c0nm_b0m_v0m_buffers0_2_, 
  c0nm_b0m_v0m_buffers0_3_, 
  c0nm_b0m_v0m_buffers0_4_, 
  c0nm_b0m_v0m_buffers0_5_, 
  c0nm_b0m_v0m_buffers0_6_, 
  c0nm_b0m_v0m_buffers0_7_, 
  c0nm_b0m_v0m_buffers0_8_, 
  c0nm_b0m_v0m_buffers0_9_, 
  c0nm_b0m_v0m_n113, 
  c0nm_b0m_v0m_n115, 
  c0nm_b0m_v0m_n134, 
  c0nm_b0m_v0m_n141, 
  c0nm_b0m_v0m_n147, 
  c0nm_b0m_v0m_n153, 
  c0nm_b0m_v0m_n159, 
  c0nm_b0m_v0m_n165, 
  c0nm_b0m_v0m_n171, 
  c0nm_b0m_v0m_n177, 
  c0nm_b0m_v0m_n183, 
  c0nm_b0m_v0m_n190, 
  c0nm_b0m_v0m_n133,
  c0nm_b0m_v0m_n140,
  c0nm_b0m_v0m_n146,
  c0nm_b0m_v0m_n152,
  c0nm_b0m_v0m_n158,
  c0nm_b0m_v0m_n164,
  c0nm_b0m_v0m_n170,
  c0nm_b0m_v0m_n176,
  c0nm_b0m_v0m_n182,
  c0nm_b0m_v0m_n189
);
  input c0nm_b0m_v0m_buffers0_10_;
  input c0nm_b0m_v0m_buffers0_11_;
  input c0nm_b0m_v0m_buffers0_2_;
  input c0nm_b0m_v0m_buffers0_3_;
  input c0nm_b0m_v0m_buffers0_4_;
  input c0nm_b0m_v0m_buffers0_5_;
  input c0nm_b0m_v0m_buffers0_6_;
  input c0nm_b0m_v0m_buffers0_7_;
  input c0nm_b0m_v0m_buffers0_8_;
  input c0nm_b0m_v0m_buffers0_9_;
  input c0nm_b0m_v0m_n113;
  input c0nm_b0m_v0m_n115;
  input c0nm_b0m_v0m_n134;
  input c0nm_b0m_v0m_n141;
  input c0nm_b0m_v0m_n147;
  input c0nm_b0m_v0m_n153;
  input c0nm_b0m_v0m_n159;
  input c0nm_b0m_v0m_n165;
  input c0nm_b0m_v0m_n171;
  input c0nm_b0m_v0m_n177;
  input c0nm_b0m_v0m_n183;
  input c0nm_b0m_v0m_n190;
  output c0nm_b0m_v0m_n133;
  output c0nm_b0m_v0m_n140;
  output c0nm_b0m_v0m_n146;
  output c0nm_b0m_v0m_n152;
  output c0nm_b0m_v0m_n158;
  output c0nm_b0m_v0m_n164;
  output c0nm_b0m_v0m_n170;
  output c0nm_b0m_v0m_n176;
  output c0nm_b0m_v0m_n182;
  output c0nm_b0m_v0m_n189;

  // moduleNum: x16
  // type: mux21i_aoi22
  // conflicting modules: 
  // number of bit inputs: 22
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 271/281
  // type: INFERRED
  // marked bad? no
  // output word of size 10 : index:99 c0nm_b0m_v0m_n170 c0nm_b0m_v0m_n146 c0nm_b0m_v0m_n133 c0nm_b0m_v0m_n140
  // c0nm_b0m_v0m_n152 c0nm_b0m_v0m_n164 c0nm_b0m_v0m_n158 c0nm_b0m_v0m_n189 c0nm_b0m_v0m_n182 c0nm_b0m_v0m_n176
  // group: sel; nodes: [ c0nm_b0m_v0m_n115 c0nm_b0m_v0m_n113 ]

  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u170 (.A0(c0nm_b0m_v0m_n115), .A1(c0nm_b0m_v0m_buffers0_11_), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n190), .Y(c0nm_b0m_v0m_n189));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u158 (.A0(c0nm_b0m_v0m_buffers0_10_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n183), .Y(c0nm_b0m_v0m_n182));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u151 (.A0(c0nm_b0m_v0m_buffers0_9_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n177), .Y(c0nm_b0m_v0m_n176));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u144 (.A0(c0nm_b0m_v0m_buffers0_8_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n171), .Y(c0nm_b0m_v0m_n170));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u137 (.A0(c0nm_b0m_v0m_buffers0_7_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n165), .Y(c0nm_b0m_v0m_n164));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u130 (.A0(c0nm_b0m_v0m_buffers0_6_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n159), .Y(c0nm_b0m_v0m_n158));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u123 (.A0(c0nm_b0m_v0m_buffers0_5_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n153), .Y(c0nm_b0m_v0m_n152));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u116 (.A0(c0nm_b0m_v0m_buffers0_4_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n147), .Y(c0nm_b0m_v0m_n146));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u109 (.A0(c0nm_b0m_v0m_buffers0_3_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n141), .Y(c0nm_b0m_v0m_n140));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u102 (.A0(c0nm_b0m_v0m_buffers0_2_), .A1(c0nm_b0m_v0m_n115), .B0(c0nm_b0m_v0m_n113), .B1(c0nm_b0m_v0m_n134), .Y(c0nm_b0m_v0m_n133));
endmodule
module mux21i_aoi22_mx17 
(
  c0sm_b0m_n2, 
  c0sm_b0m_v0m_n114, 
  c0sm_b0m_v0m_n119, 
  c0sm_b0m_v0m_n125, 
  flitin_1_0_, 
  flitin_1_1_, 
  c0sm_b0m_v0m_n118,
  c0sm_b0m_v0m_n127
);
  input c0sm_b0m_n2;
  input c0sm_b0m_v0m_n114;
  input c0sm_b0m_v0m_n119;
  input c0sm_b0m_v0m_n125;
  input flitin_1_0_;
  input flitin_1_1_;
  output c0sm_b0m_v0m_n118;
  output c0sm_b0m_v0m_n127;

  // moduleNum: x17
  // type: mux21i_aoi22
  // conflicting modules: 
  // number of bit inputs: 6
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 282/282
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:100 c0sm_b0m_v0m_n127 c0sm_b0m_v0m_n118 
  // group: sel; nodes: [ c0sm_b0m_n2 c0sm_b0m_v0m_n119 ]

  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u96 (.A0(c0sm_b0m_v0m_n119), .A1(c0sm_b0m_v0m_n125), .B0(flitin_1_1_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n127));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u89 (.A0(c0sm_b0m_v0m_n119), .A1(c0sm_b0m_v0m_n114), .B0(flitin_1_0_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n118));
endmodule
module mux21i_aoi22_mx18 
(
  c0sm_b0m_n2, 
  c0sm_b0m_v0m_buffers3_10_, 
  c0sm_b0m_v0m_buffers3_11_, 
  c0sm_b0m_v0m_buffers3_2_, 
  c0sm_b0m_v0m_buffers3_3_, 
  c0sm_b0m_v0m_buffers3_4_, 
  c0sm_b0m_v0m_buffers3_5_, 
  c0sm_b0m_v0m_buffers3_6_, 
  c0sm_b0m_v0m_buffers3_7_, 
  c0sm_b0m_v0m_buffers3_8_, 
  c0sm_b0m_v0m_buffers3_9_, 
  c0sm_b0m_v0m_n128, 
  c0sm_b0m_wdata_10_, 
  c0sm_b0m_wdata_11_, 
  c0sm_b0m_wdata_2_, 
  c0sm_b0m_wdata_3_, 
  c0sm_b0m_wdata_4_, 
  c0sm_b0m_wdata_5_, 
  c0sm_b0m_wdata_6_, 
  c0sm_b0m_wdata_7_, 
  c0sm_b0m_wdata_8_, 
  c0sm_b0m_wdata_9_, 
  flitin_1_10_, 
  flitin_1_11_, 
  flitin_1_2_, 
  flitin_1_3_, 
  flitin_1_4_, 
  flitin_1_5_, 
  flitin_1_6_, 
  flitin_1_7_, 
  flitin_1_8_, 
  flitin_1_9_, 
  c0sm_b0m_v0m_n137,
  c0sm_b0m_v0m_n143,
  c0sm_b0m_v0m_n149,
  c0sm_b0m_v0m_n155,
  c0sm_b0m_v0m_n161,
  c0sm_b0m_v0m_n167,
  c0sm_b0m_v0m_n173,
  c0sm_b0m_v0m_n179,
  c0sm_b0m_v0m_n185,
  c0sm_b0m_v0m_n195
);
  input c0sm_b0m_n2;
  input c0sm_b0m_v0m_buffers3_10_;
  input c0sm_b0m_v0m_buffers3_11_;
  input c0sm_b0m_v0m_buffers3_2_;
  input c0sm_b0m_v0m_buffers3_3_;
  input c0sm_b0m_v0m_buffers3_4_;
  input c0sm_b0m_v0m_buffers3_5_;
  input c0sm_b0m_v0m_buffers3_6_;
  input c0sm_b0m_v0m_buffers3_7_;
  input c0sm_b0m_v0m_buffers3_8_;
  input c0sm_b0m_v0m_buffers3_9_;
  input c0sm_b0m_v0m_n128;
  input c0sm_b0m_wdata_10_;
  input c0sm_b0m_wdata_11_;
  input c0sm_b0m_wdata_2_;
  input c0sm_b0m_wdata_3_;
  input c0sm_b0m_wdata_4_;
  input c0sm_b0m_wdata_5_;
  input c0sm_b0m_wdata_6_;
  input c0sm_b0m_wdata_7_;
  input c0sm_b0m_wdata_8_;
  input c0sm_b0m_wdata_9_;
  input flitin_1_10_;
  input flitin_1_11_;
  input flitin_1_2_;
  input flitin_1_3_;
  input flitin_1_4_;
  input flitin_1_5_;
  input flitin_1_6_;
  input flitin_1_7_;
  input flitin_1_8_;
  input flitin_1_9_;
  output c0sm_b0m_v0m_n137;
  output c0sm_b0m_v0m_n143;
  output c0sm_b0m_v0m_n149;
  output c0sm_b0m_v0m_n155;
  output c0sm_b0m_v0m_n161;
  output c0sm_b0m_v0m_n167;
  output c0sm_b0m_v0m_n173;
  output c0sm_b0m_v0m_n179;
  output c0sm_b0m_v0m_n185;
  output c0sm_b0m_v0m_n195;

  // moduleNum: x18
  // type: mux21i_aoi22
  // conflicting modules: 
  // number of bit inputs: 32
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 283/303
  // type: INFERRED
  // marked bad? no
  // output word of size 20 : index:101 c0sm_b0m_v0m_n143 c0sm_b0m_v0m_n143 c0sm_b0m_v0m_n137 c0sm_b0m_v0m_n137
  // c0sm_b0m_v0m_n149 c0sm_b0m_v0m_n149 c0sm_b0m_v0m_n195 c0sm_b0m_v0m_n195 c0sm_b0m_v0m_n185 c0sm_b0m_v0m_n185
  // c0sm_b0m_v0m_n179 c0sm_b0m_v0m_n179 c0sm_b0m_v0m_n173 c0sm_b0m_v0m_n173 c0sm_b0m_v0m_n167 c0sm_b0m_v0m_n167
  // c0sm_b0m_v0m_n161 c0sm_b0m_v0m_n161 c0sm_b0m_v0m_n155 c0sm_b0m_v0m_n155
  // group: sel; nodes: [ c0sm_b0m_n2 c0sm_b0m_v0m_n128 ]

  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u181 (.A0(c0sm_b0m_v0m_buffers3_11_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_n2), .B1(c0sm_b0m_wdata_11_), .Y(c0sm_b0m_v0m_n195));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u160 (.A0(c0sm_b0m_v0m_buffers3_10_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_10_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n185));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u153 (.A0(c0sm_b0m_v0m_buffers3_9_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_9_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n179));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u146 (.A0(c0sm_b0m_v0m_buffers3_8_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_8_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n173));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u139 (.A0(c0sm_b0m_v0m_buffers3_7_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_7_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n167));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u132 (.A0(c0sm_b0m_v0m_buffers3_6_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_6_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n161));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u125 (.A0(c0sm_b0m_v0m_buffers3_5_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_5_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n155));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u118 (.A0(c0sm_b0m_v0m_buffers3_4_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_4_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n149));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u111 (.A0(c0sm_b0m_v0m_buffers3_3_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_3_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n143));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u104 (.A0(c0sm_b0m_v0m_buffers3_2_), .A1(c0sm_b0m_v0m_n128), .B0(c0sm_b0m_wdata_2_), .B1(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n137));
endmodule
module mux21i_aoi22_mx19 
(
  c0sm_b0m_v0m_buffers0_3_, 
  c0sm_b0m_v0m_buffers0_5_, 
  c0sm_b0m_v0m_buffers0_6_, 
  c0sm_b0m_v0m_n141, 
  c0sm_b0m_v0m_n153, 
  c0sm_b0m_v0m_n159, 
  c0sm_b0m_v0m_n192, 
  c0sm_b0m_v0m_n193, 
  c0sm_b0m_v0m_n268,
  c0sm_b0m_v0m_n269,
  c0sm_b0m_v0m_n271
);
  input c0sm_b0m_v0m_buffers0_3_;
  input c0sm_b0m_v0m_buffers0_5_;
  input c0sm_b0m_v0m_buffers0_6_;
  input c0sm_b0m_v0m_n141;
  input c0sm_b0m_v0m_n153;
  input c0sm_b0m_v0m_n159;
  input c0sm_b0m_v0m_n192;
  input c0sm_b0m_v0m_n193;
  output c0sm_b0m_v0m_n268;
  output c0sm_b0m_v0m_n269;
  output c0sm_b0m_v0m_n271;

  // moduleNum: x19
  // type: mux21i_aoi22
  // conflicting modules: 
  // number of bit inputs: 8
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 3
  // number of non-inferred gates: 0
  // ILP vars: 334/346
  // type: INFERRED
  // marked bad? no
  // output word of size 3 : index:241 c0sm_b0m_v0m_n271 c0sm_b0m_v0m_n269 c0sm_b0m_v0m_n268 
  // group: sel; nodes: [ c0sm_b0m_v0m_n193 c0sm_b0m_v0m_n192 ]

  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u241 (.A0(c0sm_b0m_v0m_buffers0_3_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n141), .Y(c0sm_b0m_v0m_n271));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u231 (.A0(c0sm_b0m_v0m_buffers0_5_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n153), .Y(c0sm_b0m_v0m_n269));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u226 (.A0(c0sm_b0m_v0m_buffers0_6_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n159), .Y(c0sm_b0m_v0m_n268));
endmodule
module mux21i_aoi22_mx20 
(
  c0sm_b0m_v0m_buffers0_0_, 
  c0sm_b0m_v0m_buffers0_10_, 
  c0sm_b0m_v0m_buffers0_11_, 
  c0sm_b0m_v0m_buffers0_1_, 
  c0sm_b0m_v0m_buffers0_2_, 
  c0sm_b0m_v0m_buffers0_3_, 
  c0sm_b0m_v0m_buffers0_4_, 
  c0sm_b0m_v0m_buffers0_5_, 
  c0sm_b0m_v0m_buffers0_6_, 
  c0sm_b0m_v0m_buffers0_7_, 
  c0sm_b0m_v0m_buffers0_8_, 
  c0sm_b0m_v0m_buffers0_9_, 
  c0sm_b0m_v0m_buffers2_0_, 
  c0sm_b0m_v0m_buffers2_10_, 
  c0sm_b0m_v0m_buffers2_11_, 
  c0sm_b0m_v0m_buffers2_1_, 
  c0sm_b0m_v0m_buffers2_2_, 
  c0sm_b0m_v0m_buffers2_3_, 
  c0sm_b0m_v0m_buffers2_4_, 
  c0sm_b0m_v0m_buffers2_5_, 
  c0sm_b0m_v0m_buffers2_6_, 
  c0sm_b0m_v0m_buffers2_7_, 
  c0sm_b0m_v0m_buffers2_8_, 
  c0sm_b0m_v0m_buffers2_9_, 
  c0sm_b0m_v0m_n120, 
  c0sm_b0m_v0m_n121, 
  c0sm_b0m_v0m_n117,
  c0sm_b0m_v0m_n126,
  c0sm_b0m_v0m_n136,
  c0sm_b0m_v0m_n142,
  c0sm_b0m_v0m_n148,
  c0sm_b0m_v0m_n154,
  c0sm_b0m_v0m_n160,
  c0sm_b0m_v0m_n166,
  c0sm_b0m_v0m_n172,
  c0sm_b0m_v0m_n178,
  c0sm_b0m_v0m_n184,
  c0sm_b0m_v0m_n194
);
  input c0sm_b0m_v0m_buffers0_0_;
  input c0sm_b0m_v0m_buffers0_10_;
  input c0sm_b0m_v0m_buffers0_11_;
  input c0sm_b0m_v0m_buffers0_1_;
  input c0sm_b0m_v0m_buffers0_2_;
  input c0sm_b0m_v0m_buffers0_3_;
  input c0sm_b0m_v0m_buffers0_4_;
  input c0sm_b0m_v0m_buffers0_5_;
  input c0sm_b0m_v0m_buffers0_6_;
  input c0sm_b0m_v0m_buffers0_7_;
  input c0sm_b0m_v0m_buffers0_8_;
  input c0sm_b0m_v0m_buffers0_9_;
  input c0sm_b0m_v0m_buffers2_0_;
  input c0sm_b0m_v0m_buffers2_10_;
  input c0sm_b0m_v0m_buffers2_11_;
  input c0sm_b0m_v0m_buffers2_1_;
  input c0sm_b0m_v0m_buffers2_2_;
  input c0sm_b0m_v0m_buffers2_3_;
  input c0sm_b0m_v0m_buffers2_4_;
  input c0sm_b0m_v0m_buffers2_5_;
  input c0sm_b0m_v0m_buffers2_6_;
  input c0sm_b0m_v0m_buffers2_7_;
  input c0sm_b0m_v0m_buffers2_8_;
  input c0sm_b0m_v0m_buffers2_9_;
  input c0sm_b0m_v0m_n120;
  input c0sm_b0m_v0m_n121;
  output c0sm_b0m_v0m_n117;
  output c0sm_b0m_v0m_n126;
  output c0sm_b0m_v0m_n136;
  output c0sm_b0m_v0m_n142;
  output c0sm_b0m_v0m_n148;
  output c0sm_b0m_v0m_n154;
  output c0sm_b0m_v0m_n160;
  output c0sm_b0m_v0m_n166;
  output c0sm_b0m_v0m_n172;
  output c0sm_b0m_v0m_n178;
  output c0sm_b0m_v0m_n184;
  output c0sm_b0m_v0m_n194;

  // moduleNum: x20
  // type: mux21i_aoi22
  // conflicting modules: 
  // number of bit inputs: 26
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 12
  // number of non-inferred gates: 0
  // ILP vars: 377/389
  // type: INFERRED
  // marked bad? no
  // output word of size 12 : index:123 c0sm_b0m_v0m_n184 c0sm_b0m_v0m_n194 c0sm_b0m_v0m_n142 c0sm_b0m_v0m_n136
  // c0sm_b0m_v0m_n126 c0sm_b0m_v0m_n117 c0sm_b0m_v0m_n178 c0sm_b0m_v0m_n172 c0sm_b0m_v0m_n166 c0sm_b0m_v0m_n160
  // c0sm_b0m_v0m_n154 c0sm_b0m_v0m_n148
  // group: sel; nodes: [ c0sm_b0m_v0m_n121 c0sm_b0m_v0m_n120 ]

  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u184 (.A0(c0sm_b0m_v0m_buffers2_11_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_11_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n194));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u161 (.A0(c0sm_b0m_v0m_buffers2_10_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_10_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n184));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u154 (.A0(c0sm_b0m_v0m_buffers2_9_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_9_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n178));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u147 (.A0(c0sm_b0m_v0m_buffers2_8_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_8_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n172));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u140 (.A0(c0sm_b0m_v0m_buffers2_7_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_7_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n166));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u133 (.A0(c0sm_b0m_v0m_buffers2_6_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_6_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n160));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u126 (.A0(c0sm_b0m_v0m_buffers2_5_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_5_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n154));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u119 (.A0(c0sm_b0m_v0m_buffers2_4_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_4_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n148));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u112 (.A0(c0sm_b0m_v0m_buffers2_3_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_3_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n142));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u105 (.A0(c0sm_b0m_v0m_buffers2_2_), .A1(c0sm_b0m_v0m_n121), .B0(c0sm_b0m_v0m_buffers0_2_), .B1(c0sm_b0m_v0m_n120), .Y(c0sm_b0m_v0m_n136));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u97 (.A0(c0sm_b0m_v0m_buffers0_1_), .A1(c0sm_b0m_v0m_n120), .B0(c0sm_b0m_v0m_buffers2_1_), .B1(c0sm_b0m_v0m_n121), .Y(c0sm_b0m_v0m_n126));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u90 (.A0(c0sm_b0m_v0m_buffers0_0_), .A1(c0sm_b0m_v0m_n120), .B0(c0sm_b0m_v0m_buffers2_0_), .B1(c0sm_b0m_v0m_n121), .Y(c0sm_b0m_v0m_n117));
endmodule
module mux21i_aoi22_mx21 
(
  c0sm_b0m_v0m_buffers0_10_, 
  c0sm_b0m_v0m_buffers0_11_, 
  c0sm_b0m_v0m_buffers0_2_, 
  c0sm_b0m_v0m_buffers0_3_, 
  c0sm_b0m_v0m_buffers0_4_, 
  c0sm_b0m_v0m_buffers0_5_, 
  c0sm_b0m_v0m_buffers0_6_, 
  c0sm_b0m_v0m_buffers0_7_, 
  c0sm_b0m_v0m_buffers0_8_, 
  c0sm_b0m_v0m_buffers0_9_, 
  c0sm_b0m_v0m_n113, 
  c0sm_b0m_v0m_n115, 
  c0sm_b0m_v0m_n134, 
  c0sm_b0m_v0m_n141, 
  c0sm_b0m_v0m_n147, 
  c0sm_b0m_v0m_n153, 
  c0sm_b0m_v0m_n159, 
  c0sm_b0m_v0m_n165, 
  c0sm_b0m_v0m_n171, 
  c0sm_b0m_v0m_n177, 
  c0sm_b0m_v0m_n183, 
  c0sm_b0m_v0m_n190, 
  c0sm_b0m_v0m_n133,
  c0sm_b0m_v0m_n140,
  c0sm_b0m_v0m_n146,
  c0sm_b0m_v0m_n152,
  c0sm_b0m_v0m_n158,
  c0sm_b0m_v0m_n164,
  c0sm_b0m_v0m_n170,
  c0sm_b0m_v0m_n176,
  c0sm_b0m_v0m_n182,
  c0sm_b0m_v0m_n189
);
  input c0sm_b0m_v0m_buffers0_10_;
  input c0sm_b0m_v0m_buffers0_11_;
  input c0sm_b0m_v0m_buffers0_2_;
  input c0sm_b0m_v0m_buffers0_3_;
  input c0sm_b0m_v0m_buffers0_4_;
  input c0sm_b0m_v0m_buffers0_5_;
  input c0sm_b0m_v0m_buffers0_6_;
  input c0sm_b0m_v0m_buffers0_7_;
  input c0sm_b0m_v0m_buffers0_8_;
  input c0sm_b0m_v0m_buffers0_9_;
  input c0sm_b0m_v0m_n113;
  input c0sm_b0m_v0m_n115;
  input c0sm_b0m_v0m_n134;
  input c0sm_b0m_v0m_n141;
  input c0sm_b0m_v0m_n147;
  input c0sm_b0m_v0m_n153;
  input c0sm_b0m_v0m_n159;
  input c0sm_b0m_v0m_n165;
  input c0sm_b0m_v0m_n171;
  input c0sm_b0m_v0m_n177;
  input c0sm_b0m_v0m_n183;
  input c0sm_b0m_v0m_n190;
  output c0sm_b0m_v0m_n133;
  output c0sm_b0m_v0m_n140;
  output c0sm_b0m_v0m_n146;
  output c0sm_b0m_v0m_n152;
  output c0sm_b0m_v0m_n158;
  output c0sm_b0m_v0m_n164;
  output c0sm_b0m_v0m_n170;
  output c0sm_b0m_v0m_n176;
  output c0sm_b0m_v0m_n182;
  output c0sm_b0m_v0m_n189;

  // moduleNum: x21
  // type: mux21i_aoi22
  // conflicting modules: 
  // number of bit inputs: 22
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 420/430
  // type: INFERRED
  // marked bad? no
  // output word of size 10 : index:124 c0sm_b0m_v0m_n170 c0sm_b0m_v0m_n133 c0sm_b0m_v0m_n164 c0sm_b0m_v0m_n140
  // c0sm_b0m_v0m_n158 c0sm_b0m_v0m_n146 c0sm_b0m_v0m_n152 c0sm_b0m_v0m_n189 c0sm_b0m_v0m_n182 c0sm_b0m_v0m_n176
  // group: sel; nodes: [ c0sm_b0m_v0m_n115 c0sm_b0m_v0m_n113 ]

  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u170 (.A0(c0sm_b0m_v0m_n115), .A1(c0sm_b0m_v0m_buffers0_11_), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n190), .Y(c0sm_b0m_v0m_n189));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u158 (.A0(c0sm_b0m_v0m_buffers0_10_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n183), .Y(c0sm_b0m_v0m_n182));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u151 (.A0(c0sm_b0m_v0m_buffers0_9_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n177), .Y(c0sm_b0m_v0m_n176));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u144 (.A0(c0sm_b0m_v0m_buffers0_8_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n171), .Y(c0sm_b0m_v0m_n170));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u137 (.A0(c0sm_b0m_v0m_buffers0_7_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n165), .Y(c0sm_b0m_v0m_n164));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u130 (.A0(c0sm_b0m_v0m_buffers0_6_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n159), .Y(c0sm_b0m_v0m_n158));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u123 (.A0(c0sm_b0m_v0m_buffers0_5_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n153), .Y(c0sm_b0m_v0m_n152));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u116 (.A0(c0sm_b0m_v0m_buffers0_4_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n147), .Y(c0sm_b0m_v0m_n146));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u109 (.A0(c0sm_b0m_v0m_buffers0_3_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n141), .Y(c0sm_b0m_v0m_n140));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u102 (.A0(c0sm_b0m_v0m_buffers0_2_), .A1(c0sm_b0m_v0m_n115), .B0(c0sm_b0m_v0m_n113), .B1(c0sm_b0m_v0m_n134), .Y(c0sm_b0m_v0m_n133));
endmodule
module mux31b_mx22 
(
  flitout_switch_0_0_, 
  flitout_switch_0_10_, 
  flitout_switch_0_11_, 
  flitout_switch_0_1_, 
  flitout_switch_0_2_, 
  flitout_switch_0_3_, 
  flitout_switch_0_4_, 
  flitout_switch_0_5_, 
  flitout_switch_0_6_, 
  flitout_switch_0_7_, 
  flitout_switch_0_8_, 
  flitout_switch_0_9_, 
  flitout_switch_1_0_, 
  flitout_switch_1_10_, 
  flitout_switch_1_11_, 
  flitout_switch_1_1_, 
  flitout_switch_1_2_, 
  flitout_switch_1_3_, 
  flitout_switch_1_4_, 
  flitout_switch_1_5_, 
  flitout_switch_1_6_, 
  flitout_switch_1_7_, 
  flitout_switch_1_8_, 
  flitout_switch_1_9_, 
  x0m__logic0_, 
  x0m__logic1_, 
  x0m_colsel0reg_0_, 
  x0m_colsel0reg_1_, 
  flitout_0_0_,
  flitout_0_10_,
  flitout_0_11_,
  flitout_0_1_,
  flitout_0_2_,
  flitout_0_3_,
  flitout_0_4_,
  flitout_0_5_,
  flitout_0_6_,
  flitout_0_7_,
  flitout_0_8_,
  flitout_0_9_
);
  input flitout_switch_0_0_;
  input flitout_switch_0_10_;
  input flitout_switch_0_11_;
  input flitout_switch_0_1_;
  input flitout_switch_0_2_;
  input flitout_switch_0_3_;
  input flitout_switch_0_4_;
  input flitout_switch_0_5_;
  input flitout_switch_0_6_;
  input flitout_switch_0_7_;
  input flitout_switch_0_8_;
  input flitout_switch_0_9_;
  input flitout_switch_1_0_;
  input flitout_switch_1_10_;
  input flitout_switch_1_11_;
  input flitout_switch_1_1_;
  input flitout_switch_1_2_;
  input flitout_switch_1_3_;
  input flitout_switch_1_4_;
  input flitout_switch_1_5_;
  input flitout_switch_1_6_;
  input flitout_switch_1_7_;
  input flitout_switch_1_8_;
  input flitout_switch_1_9_;
  input x0m__logic0_;
  input x0m__logic1_;
  input x0m_colsel0reg_0_;
  input x0m_colsel0reg_1_;
  output flitout_0_0_;
  output flitout_0_10_;
  output flitout_0_11_;
  output flitout_0_1_;
  output flitout_0_2_;
  output flitout_0_3_;
  output flitout_0_4_;
  output flitout_0_5_;
  output flitout_0_6_;
  output flitout_0_7_;
  output flitout_0_8_;
  output flitout_0_9_;
  wire x0m_bx0m_m0m_int01;
  wire x0m_bx10m_m0m_int01;
  wire x0m_bx11m_m0m_int01;
  wire x0m_bx1m_m0m_int01;
  wire x0m_bx2m_m0m_int01;
  wire x0m_bx3m_m0m_int01;
  wire x0m_bx4m_m0m_int01;
  wire x0m_bx5m_m0m_int01;
  wire x0m_bx6m_m0m_int01;
  wire x0m_bx7m_m0m_int01;
  wire x0m_bx8m_m0m_int01;
  wire x0m_bx9m_m0m_int01;

  // moduleNum: x22
  // type: mux31b
  // conflicting modules: 
  // number of bit inputs: 2
  // number of bit outputs: 0
  // number of word inputs: 3
  // number of word outputs: 1
  // number of internal gates: 24
  // number of non-inferred gates: 0
  // ILP vars: 431/443
  // type: INFERRED
  // marked bad? no
  // input word of size 12 : index:125 flitout_switch_0[6] flitout_switch_0[5] flitout_switch_0[4] flitout_switch_0[3]
  // flitout_switch_0[2] flitout_switch_0[1] flitout_switch_0[11] flitout_switch_0[0] flitout_switch_0[10]
  // flitout_switch_0[7] flitout_switch_0[8] flitout_switch_0[9]
  // input word of size 12 : index:126 flitout_switch_1[6] flitout_switch_1[5] flitout_switch_1[4] flitout_switch_1[3]
  // flitout_switch_1[2] flitout_switch_1[1] flitout_switch_1[11] flitout_switch_1[0] flitout_switch_1[10]
  // flitout_switch_1[7] flitout_switch_1[8] flitout_switch_1[9]
  // input word of size 12 : index:16 x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic1_
  // x0m__logic0_ x0m__logic1_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_
  // output word of size 12 : index:17 flitout_0[6] flitout_0[5] flitout_0[4] flitout_0[3] flitout_0[2] flitout_0[1]
  // flitout_0[11] flitout_0[0] flitout_0[10] flitout_0[7] flitout_0[8] flitout_0[9]
  // group: sel; nodes: [ x0m_colsel0reg_0_ x0m_colsel0reg_1_ ]

  MXT2_X0P5M_A12TR x0m_bx0m_m0m_m0m_u1 (.A(flitout_switch_0_0_), .B(flitout_switch_1_0_), .S0(x0m_colsel0reg_0_), .Y(x0m_bx0m_m0m_int01));
  MXT2_X0P5M_A12TR x0m_bx0m_m0m_m4m_u1 (.A(x0m_bx0m_m0m_int01), .B(x0m__logic1_), .S0(x0m_colsel0reg_1_), .Y(flitout_0_0_));
  MXT2_X0P5M_A12TR x0m_bx1m_m0m_m0m_u1 (.A(flitout_switch_0_1_), .B(flitout_switch_1_1_), .S0(x0m_colsel0reg_0_), .Y(x0m_bx1m_m0m_int01));
  MXT2_X0P5M_A12TR x0m_bx1m_m0m_m4m_u1 (.A(x0m_bx1m_m0m_int01), .B(x0m__logic1_), .S0(x0m_colsel0reg_1_), .Y(flitout_0_1_));
  MXT2_X0P5M_A12TR x0m_bx2m_m0m_m0m_u1 (.A(flitout_switch_0_2_), .B(flitout_switch_1_2_), .S0(x0m_colsel0reg_0_), .Y(x0m_bx2m_m0m_int01));
  MXT2_X0P5M_A12TR x0m_bx2m_m0m_m4m_u1 (.A(x0m_bx2m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0_2_));
  MXT2_X0P5M_A12TR x0m_bx3m_m0m_m0m_u1 (.A(flitout_switch_0_3_), .B(flitout_switch_1_3_), .S0(x0m_colsel0reg_0_), .Y(x0m_bx3m_m0m_int01));
  MXT2_X0P5M_A12TR x0m_bx3m_m0m_m4m_u1 (.A(x0m_bx3m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0_3_));
  MXT2_X0P5M_A12TR x0m_bx4m_m0m_m0m_u1 (.A(flitout_switch_0_4_), .B(flitout_switch_1_4_), .S0(x0m_colsel0reg_0_), .Y(x0m_bx4m_m0m_int01));
  MXT2_X0P5M_A12TR x0m_bx4m_m0m_m4m_u1 (.A(x0m_bx4m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0_4_));
  MXT2_X0P5M_A12TR x0m_bx5m_m0m_m0m_u1 (.A(flitout_switch_0_5_), .B(flitout_switch_1_5_), .S0(x0m_colsel0reg_0_), .Y(x0m_bx5m_m0m_int01));
  MXT2_X0P5M_A12TR x0m_bx5m_m0m_m4m_u1 (.A(x0m_bx5m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0_5_));
  MXT2_X0P5M_A12TR x0m_bx6m_m0m_m0m_u1 (.A(flitout_switch_0_6_), .B(flitout_switch_1_6_), .S0(x0m_colsel0reg_0_), .Y(x0m_bx6m_m0m_int01));
  MXT2_X0P5M_A12TR x0m_bx6m_m0m_m4m_u1 (.A(x0m_bx6m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0_6_));
  MXT2_X0P5M_A12TR x0m_bx7m_m0m_m0m_u1 (.A(flitout_switch_0_7_), .B(flitout_switch_1_7_), .S0(x0m_colsel0reg_0_), .Y(x0m_bx7m_m0m_int01));
  MXT2_X0P5M_A12TR x0m_bx7m_m0m_m4m_u1 (.A(x0m_bx7m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0_7_));
  MXT2_X0P5M_A12TR x0m_bx8m_m0m_m0m_u1 (.A(flitout_switch_0_8_), .B(flitout_switch_1_8_), .S0(x0m_colsel0reg_0_), .Y(x0m_bx8m_m0m_int01));
  MXT2_X0P5M_A12TR x0m_bx8m_m0m_m4m_u1 (.A(x0m_bx8m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0_8_));
  MXT2_X0P5M_A12TR x0m_bx9m_m0m_m0m_u1 (.A(flitout_switch_0_9_), .B(flitout_switch_1_9_), .S0(x0m_colsel0reg_0_), .Y(x0m_bx9m_m0m_int01));
  MXT2_X0P5M_A12TR x0m_bx9m_m0m_m4m_u1 (.A(x0m_bx9m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0_9_));
  MXT2_X0P5M_A12TR x0m_bx10m_m0m_m0m_u1 (.A(flitout_switch_0_10_), .B(flitout_switch_1_10_), .S0(x0m_colsel0reg_0_), .Y(x0m_bx10m_m0m_int01));
  MXT2_X0P5M_A12TR x0m_bx10m_m0m_m4m_u1 (.A(x0m_bx10m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0_10_));
  MXT2_X0P5M_A12TR x0m_bx11m_m0m_m0m_u1 (.A(flitout_switch_0_11_), .B(flitout_switch_1_11_), .S0(x0m_colsel0reg_0_), .Y(x0m_bx11m_m0m_int01));
  MXT2_X0P5M_A12TR x0m_bx11m_m0m_m4m_u1 (.A(x0m_bx11m_m0m_int01), .B(x0m__logic0_), .S0(x0m_colsel0reg_1_), .Y(flitout_0_11_));
endmodule
module mux31b_mx23 
(
  flitout_switch_0_10_, 
  flitout_switch_0_2_, 
  flitout_switch_0_3_, 
  flitout_switch_0_5_, 
  flitout_switch_0_6_, 
  flitout_switch_0_7_, 
  flitout_switch_0_8_, 
  flitout_switch_0_9_, 
  flitout_switch_1_10_, 
  flitout_switch_1_2_, 
  flitout_switch_1_3_, 
  flitout_switch_1_5_, 
  flitout_switch_1_6_, 
  flitout_switch_1_7_, 
  flitout_switch_1_8_, 
  flitout_switch_1_9_, 
  x0m__logic0_, 
  x0m_colsel1reg_0_, 
  x0m_colsel1reg_1_, 
  flitout_1_10_,
  flitout_1_2_,
  flitout_1_3_,
  flitout_1_5_,
  flitout_1_6_,
  flitout_1_7_,
  flitout_1_8_,
  flitout_1_9_
);
  input flitout_switch_0_10_;
  input flitout_switch_0_2_;
  input flitout_switch_0_3_;
  input flitout_switch_0_5_;
  input flitout_switch_0_6_;
  input flitout_switch_0_7_;
  input flitout_switch_0_8_;
  input flitout_switch_0_9_;
  input flitout_switch_1_10_;
  input flitout_switch_1_2_;
  input flitout_switch_1_3_;
  input flitout_switch_1_5_;
  input flitout_switch_1_6_;
  input flitout_switch_1_7_;
  input flitout_switch_1_8_;
  input flitout_switch_1_9_;
  input x0m__logic0_;
  input x0m_colsel1reg_0_;
  input x0m_colsel1reg_1_;
  output flitout_1_10_;
  output flitout_1_2_;
  output flitout_1_3_;
  output flitout_1_5_;
  output flitout_1_6_;
  output flitout_1_7_;
  output flitout_1_8_;
  output flitout_1_9_;
  wire x0m_bx10m_m1m_int01;
  wire x0m_bx2m_m1m_int01;
  wire x0m_bx3m_m1m_int01;
  wire x0m_bx5m_m1m_int01;
  wire x0m_bx6m_m1m_int01;
  wire x0m_bx7m_m1m_int01;
  wire x0m_bx8m_m1m_int01;
  wire x0m_bx9m_m1m_int01;

  // moduleNum: x23
  // type: mux31b
  // conflicting modules: 
  // number of bit inputs: 2
  // number of bit outputs: 0
  // number of word inputs: 3
  // number of word outputs: 1
  // number of internal gates: 16
  // number of non-inferred gates: 0
  // ILP vars: 444/455
  // type: INFERRED
  // marked bad? no
  // input word of size 8 : index:-1 flitout_switch_0[3] flitout_switch_0[2] flitout_switch_0[10] flitout_switch_0[6]
  // flitout_switch_0[7] flitout_switch_0[8] flitout_switch_0[9] flitout_switch_0[5]
  // input word of size 8 : index:-1 flitout_switch_1[3] flitout_switch_1[2] flitout_switch_1[10] flitout_switch_1[6]
  // flitout_switch_1[7] flitout_switch_1[8] flitout_switch_1[9] flitout_switch_1[5]
  // input word of size 9 : index:-1 x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_ x0m__logic0_
  // x0m__logic0_ x0m__logic0_ x0m__logic0_
  // output word of size 8 : index:242 flitout_1[3] flitout_1[2] flitout_1[10] flitout_1[6] flitout_1[7] flitout_1[8]
  // flitout_1[9] flitout_1[5]
  // group: sel; nodes: [ x0m_colsel1reg_0_ x0m_colsel1reg_1_ ]

  MXT2_X0P5M_A12TR x0m_bx2m_m1m_m0m_u1 (.A(flitout_switch_0_2_), .B(flitout_switch_1_2_), .S0(x0m_colsel1reg_0_), .Y(x0m_bx2m_m1m_int01));
  MXT2_X0P5M_A12TR x0m_bx2m_m1m_m4m_u1 (.A(x0m_bx2m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1_2_));
  MXT2_X0P5M_A12TR x0m_bx3m_m1m_m0m_u1 (.A(flitout_switch_0_3_), .B(flitout_switch_1_3_), .S0(x0m_colsel1reg_0_), .Y(x0m_bx3m_m1m_int01));
  MXT2_X0P5M_A12TR x0m_bx3m_m1m_m4m_u1 (.A(x0m_bx3m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1_3_));
  MXT2_X0P5M_A12TR x0m_bx5m_m1m_m0m_u1 (.A(flitout_switch_0_5_), .B(flitout_switch_1_5_), .S0(x0m_colsel1reg_0_), .Y(x0m_bx5m_m1m_int01));
  MXT2_X0P5M_A12TR x0m_bx5m_m1m_m4m_u1 (.A(x0m_bx5m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1_5_));
  MXT2_X0P5M_A12TR x0m_bx6m_m1m_m0m_u1 (.A(flitout_switch_0_6_), .B(flitout_switch_1_6_), .S0(x0m_colsel1reg_0_), .Y(x0m_bx6m_m1m_int01));
  MXT2_X0P5M_A12TR x0m_bx6m_m1m_m4m_u1 (.A(x0m_bx6m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1_6_));
  MXT2_X0P5M_A12TR x0m_bx7m_m1m_m0m_u1 (.A(flitout_switch_0_7_), .B(flitout_switch_1_7_), .S0(x0m_colsel1reg_0_), .Y(x0m_bx7m_m1m_int01));
  MXT2_X0P5M_A12TR x0m_bx7m_m1m_m4m_u1 (.A(x0m_bx7m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1_7_));
  MXT2_X0P5M_A12TR x0m_bx8m_m1m_m0m_u1 (.A(flitout_switch_0_8_), .B(flitout_switch_1_8_), .S0(x0m_colsel1reg_0_), .Y(x0m_bx8m_m1m_int01));
  MXT2_X0P5M_A12TR x0m_bx8m_m1m_m4m_u1 (.A(x0m_bx8m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1_8_));
  MXT2_X0P5M_A12TR x0m_bx9m_m1m_m0m_u1 (.A(flitout_switch_0_9_), .B(flitout_switch_1_9_), .S0(x0m_colsel1reg_0_), .Y(x0m_bx9m_m1m_int01));
  MXT2_X0P5M_A12TR x0m_bx9m_m1m_m4m_u1 (.A(x0m_bx9m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1_9_));
  MXT2_X0P5M_A12TR x0m_bx10m_m1m_m0m_u1 (.A(flitout_switch_0_10_), .B(flitout_switch_1_10_), .S0(x0m_colsel1reg_0_), .Y(x0m_bx10m_m1m_int01));
  MXT2_X0P5M_A12TR x0m_bx10m_m1m_m4m_u1 (.A(x0m_bx10m_m1m_int01), .B(x0m__logic0_), .S0(x0m_colsel1reg_1_), .Y(flitout_1_10_));
endmodule
module mux31i_oai222_mx24 
(
  c0nm_b0m_v0m_n107, 
  c0nm_b0m_v0m_n129, 
  c0nm_b0m_v0m_n130, 
  c0nm_b0m_v0m_n131, 
  c0nm_b0m_v0m_n138, 
  c0nm_b0m_v0m_n144, 
  c0nm_b0m_v0m_n150, 
  c0nm_b0m_v0m_n156, 
  c0nm_b0m_v0m_n162, 
  c0nm_b0m_v0m_n168, 
  c0nm_b0m_v0m_n17, 
  c0nm_b0m_v0m_n174, 
  c0nm_b0m_v0m_n180, 
  c0nm_b0m_v0m_n186, 
  c0nm_b0m_v0m_n19, 
  c0nm_b0m_v0m_n33, 
  c0nm_b0m_v0m_n34, 
  c0nm_b0m_v0m_n36, 
  c0nm_b0m_v0m_n37, 
  c0nm_b0m_v0m_n39, 
  c0nm_b0m_v0m_n40, 
  c0nm_b0m_v0m_n42, 
  c0nm_b0m_v0m_n43, 
  c0nm_b0m_v0m_n45, 
  c0nm_b0m_v0m_n46, 
  c0nm_b0m_v0m_n48, 
  c0nm_b0m_v0m_n49, 
  c0nm_b0m_v0m_n63, 
  c0nm_b0m_v0m_n64, 
  c0nm_b0m_v0m_n66, 
  c0nm_b0m_v0m_n67, 
  c0nm_b0m_v0m_n69, 
  c0nm_b0m_v0m_n70, 
  c0nm_b0m_v0m_n208,
  c0nm_b0m_v0m_n209,
  c0nm_b0m_v0m_n210,
  c0nm_b0m_v0m_n211,
  c0nm_b0m_v0m_n212,
  c0nm_b0m_v0m_n213,
  c0nm_b0m_v0m_n214,
  c0nm_b0m_v0m_n215,
  c0nm_b0m_v0m_n216,
  c0nm_b0m_v0m_n217
);
  input c0nm_b0m_v0m_n107;
  input c0nm_b0m_v0m_n129;
  input c0nm_b0m_v0m_n130;
  input c0nm_b0m_v0m_n131;
  input c0nm_b0m_v0m_n138;
  input c0nm_b0m_v0m_n144;
  input c0nm_b0m_v0m_n150;
  input c0nm_b0m_v0m_n156;
  input c0nm_b0m_v0m_n162;
  input c0nm_b0m_v0m_n168;
  input c0nm_b0m_v0m_n17;
  input c0nm_b0m_v0m_n174;
  input c0nm_b0m_v0m_n180;
  input c0nm_b0m_v0m_n186;
  input c0nm_b0m_v0m_n19;
  input c0nm_b0m_v0m_n33;
  input c0nm_b0m_v0m_n34;
  input c0nm_b0m_v0m_n36;
  input c0nm_b0m_v0m_n37;
  input c0nm_b0m_v0m_n39;
  input c0nm_b0m_v0m_n40;
  input c0nm_b0m_v0m_n42;
  input c0nm_b0m_v0m_n43;
  input c0nm_b0m_v0m_n45;
  input c0nm_b0m_v0m_n46;
  input c0nm_b0m_v0m_n48;
  input c0nm_b0m_v0m_n49;
  input c0nm_b0m_v0m_n63;
  input c0nm_b0m_v0m_n64;
  input c0nm_b0m_v0m_n66;
  input c0nm_b0m_v0m_n67;
  input c0nm_b0m_v0m_n69;
  input c0nm_b0m_v0m_n70;
  output c0nm_b0m_v0m_n208;
  output c0nm_b0m_v0m_n209;
  output c0nm_b0m_v0m_n210;
  output c0nm_b0m_v0m_n211;
  output c0nm_b0m_v0m_n212;
  output c0nm_b0m_v0m_n213;
  output c0nm_b0m_v0m_n214;
  output c0nm_b0m_v0m_n215;
  output c0nm_b0m_v0m_n216;
  output c0nm_b0m_v0m_n217;

  // moduleNum: x24
  // type: mux31i_oai222
  // conflicting modules: 
  // number of bit inputs: 33
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 456/466
  // type: INFERRED
  // marked bad? no
  // output word of size 10 : index:131 c0nm_b0m_v0m_n208 c0nm_b0m_v0m_n209 c0nm_b0m_v0m_n210 c0nm_b0m_v0m_n211
  // c0nm_b0m_v0m_n212 c0nm_b0m_v0m_n213 c0nm_b0m_v0m_n214 c0nm_b0m_v0m_n215 c0nm_b0m_v0m_n216 c0nm_b0m_v0m_n217
  // group: sel; nodes: [ c0nm_b0m_v0m_n129 c0nm_b0m_v0m_n107 c0nm_b0m_v0m_n130 ]

  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u162 (.A0(c0nm_b0m_v0m_n19), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n17), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n186), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n208));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u155 (.A0(c0nm_b0m_v0m_n70), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n69), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n180), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n209));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u148 (.A0(c0nm_b0m_v0m_n67), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n66), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n174), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n210));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u141 (.A0(c0nm_b0m_v0m_n64), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n63), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n168), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n211));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u134 (.A0(c0nm_b0m_v0m_n49), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n48), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n162), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n212));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u127 (.A0(c0nm_b0m_v0m_n46), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n45), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n156), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n213));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u120 (.A0(c0nm_b0m_v0m_n43), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n42), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n150), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n214));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u113 (.A0(c0nm_b0m_v0m_n40), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n39), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n144), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n215));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u106 (.A0(c0nm_b0m_v0m_n37), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n36), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n138), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n216));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u99 (.A0(c0nm_b0m_v0m_n34), .A1(c0nm_b0m_v0m_n129), .B0(c0nm_b0m_v0m_n33), .B1(c0nm_b0m_v0m_n130), .C0(c0nm_b0m_v0m_n131), .C1(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n217));
endmodule
module mux31i_oai222_mx25 
(
  c0nm_b0m_v0m_n17, 
  c0nm_b0m_v0m_n19, 
  c0nm_b0m_v0m_n33, 
  c0nm_b0m_v0m_n34, 
  c0nm_b0m_v0m_n36, 
  c0nm_b0m_v0m_n37, 
  c0nm_b0m_v0m_n39, 
  c0nm_b0m_v0m_n40, 
  c0nm_b0m_v0m_n42, 
  c0nm_b0m_v0m_n43, 
  c0nm_b0m_v0m_n45, 
  c0nm_b0m_v0m_n46, 
  c0nm_b0m_v0m_n48, 
  c0nm_b0m_v0m_n49, 
  c0nm_b0m_v0m_n63, 
  c0nm_b0m_v0m_n64, 
  c0nm_b0m_v0m_n66, 
  c0nm_b0m_v0m_n67, 
  c0nm_b0m_v0m_n69, 
  c0nm_b0m_v0m_n70, 
  c0nm_b0m_v0m_n76, 
  c0nm_b0m_v0m_n81, 
  c0nm_b0m_v0m_n82, 
  c0nm_b0m_v0m_n83, 
  c0nm_b0m_v0m_n84, 
  c0nm_b0m_v0m_n85, 
  c0nm_b0m_v0m_n86, 
  c0nm_b0m_v0m_n87, 
  c0nm_b0m_v0m_n88, 
  c0nm_b0m_v0m_n89, 
  c0nm_b0m_v0m_n90, 
  c0nm_b0m_v0m_n91, 
  c0nm_b0m_v0m_n92, 
  c0nm_b0m_v0m_n232,
  c0nm_b0m_v0m_n233,
  c0nm_b0m_v0m_n234,
  c0nm_b0m_v0m_n235,
  c0nm_b0m_v0m_n236,
  c0nm_b0m_v0m_n237,
  c0nm_b0m_v0m_n238,
  c0nm_b0m_v0m_n239,
  c0nm_b0m_v0m_n240,
  c0nm_b0m_v0m_n241
);
  input c0nm_b0m_v0m_n17;
  input c0nm_b0m_v0m_n19;
  input c0nm_b0m_v0m_n33;
  input c0nm_b0m_v0m_n34;
  input c0nm_b0m_v0m_n36;
  input c0nm_b0m_v0m_n37;
  input c0nm_b0m_v0m_n39;
  input c0nm_b0m_v0m_n40;
  input c0nm_b0m_v0m_n42;
  input c0nm_b0m_v0m_n43;
  input c0nm_b0m_v0m_n45;
  input c0nm_b0m_v0m_n46;
  input c0nm_b0m_v0m_n48;
  input c0nm_b0m_v0m_n49;
  input c0nm_b0m_v0m_n63;
  input c0nm_b0m_v0m_n64;
  input c0nm_b0m_v0m_n66;
  input c0nm_b0m_v0m_n67;
  input c0nm_b0m_v0m_n69;
  input c0nm_b0m_v0m_n70;
  input c0nm_b0m_v0m_n76;
  input c0nm_b0m_v0m_n81;
  input c0nm_b0m_v0m_n82;
  input c0nm_b0m_v0m_n83;
  input c0nm_b0m_v0m_n84;
  input c0nm_b0m_v0m_n85;
  input c0nm_b0m_v0m_n86;
  input c0nm_b0m_v0m_n87;
  input c0nm_b0m_v0m_n88;
  input c0nm_b0m_v0m_n89;
  input c0nm_b0m_v0m_n90;
  input c0nm_b0m_v0m_n91;
  input c0nm_b0m_v0m_n92;
  output c0nm_b0m_v0m_n232;
  output c0nm_b0m_v0m_n233;
  output c0nm_b0m_v0m_n234;
  output c0nm_b0m_v0m_n235;
  output c0nm_b0m_v0m_n236;
  output c0nm_b0m_v0m_n237;
  output c0nm_b0m_v0m_n238;
  output c0nm_b0m_v0m_n239;
  output c0nm_b0m_v0m_n240;
  output c0nm_b0m_v0m_n241;

  // moduleNum: x25
  // type: mux31i_oai222
  // conflicting modules: 
  // number of bit inputs: 33
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 478/488
  // type: INFERRED
  // marked bad? no
  // output word of size 10 : index:133 c0nm_b0m_v0m_n232 c0nm_b0m_v0m_n239 c0nm_b0m_v0m_n238 c0nm_b0m_v0m_n237
  // c0nm_b0m_v0m_n236 c0nm_b0m_v0m_n235 c0nm_b0m_v0m_n234 c0nm_b0m_v0m_n233 c0nm_b0m_v0m_n241 c0nm_b0m_v0m_n240
  // group: sel; nodes: [ c0nm_b0m_v0m_n81 c0nm_b0m_v0m_n76 c0nm_b0m_v0m_n82 ]

  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u58 (.A0(c0nm_b0m_v0m_n19), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n17), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n92), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n232));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u56 (.A0(c0nm_b0m_v0m_n70), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n69), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n91), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n233));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u54 (.A0(c0nm_b0m_v0m_n67), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n66), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n90), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n234));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u52 (.A0(c0nm_b0m_v0m_n64), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n63), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n89), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n235));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u50 (.A0(c0nm_b0m_v0m_n49), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n48), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n88), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n236));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u48 (.A0(c0nm_b0m_v0m_n46), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n45), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n87), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n237));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u46 (.A0(c0nm_b0m_v0m_n43), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n42), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n86), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n238));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u44 (.A0(c0nm_b0m_v0m_n40), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n39), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n85), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n239));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u42 (.A0(c0nm_b0m_v0m_n37), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n36), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n84), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n240));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u40 (.A0(c0nm_b0m_v0m_n34), .A1(c0nm_b0m_v0m_n81), .B0(c0nm_b0m_v0m_n33), .B1(c0nm_b0m_v0m_n82), .C0(c0nm_b0m_v0m_n83), .C1(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n241));
endmodule
module mux31i_oai222_mx26 
(
  c0nm_b0m_v0m_n17, 
  c0nm_b0m_v0m_n18, 
  c0nm_b0m_v0m_n19, 
  c0nm_b0m_v0m_n20, 
  c0nm_b0m_v0m_n21, 
  c0nm_b0m_v0m_n22, 
  c0nm_b0m_v0m_n33, 
  c0nm_b0m_v0m_n34, 
  c0nm_b0m_v0m_n35, 
  c0nm_b0m_v0m_n36, 
  c0nm_b0m_v0m_n37, 
  c0nm_b0m_v0m_n38, 
  c0nm_b0m_v0m_n39, 
  c0nm_b0m_v0m_n40, 
  c0nm_b0m_v0m_n41, 
  c0nm_b0m_v0m_n42, 
  c0nm_b0m_v0m_n43, 
  c0nm_b0m_v0m_n44, 
  c0nm_b0m_v0m_n45, 
  c0nm_b0m_v0m_n46, 
  c0nm_b0m_v0m_n47, 
  c0nm_b0m_v0m_n48, 
  c0nm_b0m_v0m_n49, 
  c0nm_b0m_v0m_n62, 
  c0nm_b0m_v0m_n63, 
  c0nm_b0m_v0m_n64, 
  c0nm_b0m_v0m_n65, 
  c0nm_b0m_v0m_n66, 
  c0nm_b0m_v0m_n67, 
  c0nm_b0m_v0m_n68, 
  c0nm_b0m_v0m_n69, 
  c0nm_b0m_v0m_n70, 
  c0nm_b0m_v0m_n71, 
  c0nm_b0m_v0m_n244,
  c0nm_b0m_v0m_n245,
  c0nm_b0m_v0m_n246,
  c0nm_b0m_v0m_n247,
  c0nm_b0m_v0m_n248,
  c0nm_b0m_v0m_n249,
  c0nm_b0m_v0m_n250,
  c0nm_b0m_v0m_n251,
  c0nm_b0m_v0m_n252,
  c0nm_b0m_v0m_n255
);
  input c0nm_b0m_v0m_n17;
  input c0nm_b0m_v0m_n18;
  input c0nm_b0m_v0m_n19;
  input c0nm_b0m_v0m_n20;
  input c0nm_b0m_v0m_n21;
  input c0nm_b0m_v0m_n22;
  input c0nm_b0m_v0m_n33;
  input c0nm_b0m_v0m_n34;
  input c0nm_b0m_v0m_n35;
  input c0nm_b0m_v0m_n36;
  input c0nm_b0m_v0m_n37;
  input c0nm_b0m_v0m_n38;
  input c0nm_b0m_v0m_n39;
  input c0nm_b0m_v0m_n40;
  input c0nm_b0m_v0m_n41;
  input c0nm_b0m_v0m_n42;
  input c0nm_b0m_v0m_n43;
  input c0nm_b0m_v0m_n44;
  input c0nm_b0m_v0m_n45;
  input c0nm_b0m_v0m_n46;
  input c0nm_b0m_v0m_n47;
  input c0nm_b0m_v0m_n48;
  input c0nm_b0m_v0m_n49;
  input c0nm_b0m_v0m_n62;
  input c0nm_b0m_v0m_n63;
  input c0nm_b0m_v0m_n64;
  input c0nm_b0m_v0m_n65;
  input c0nm_b0m_v0m_n66;
  input c0nm_b0m_v0m_n67;
  input c0nm_b0m_v0m_n68;
  input c0nm_b0m_v0m_n69;
  input c0nm_b0m_v0m_n70;
  input c0nm_b0m_v0m_n71;
  output c0nm_b0m_v0m_n244;
  output c0nm_b0m_v0m_n245;
  output c0nm_b0m_v0m_n246;
  output c0nm_b0m_v0m_n247;
  output c0nm_b0m_v0m_n248;
  output c0nm_b0m_v0m_n249;
  output c0nm_b0m_v0m_n250;
  output c0nm_b0m_v0m_n251;
  output c0nm_b0m_v0m_n252;
  output c0nm_b0m_v0m_n255;

  // moduleNum: x26
  // type: mux31i_oai222
  // conflicting modules: 
  // number of bit inputs: 33
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 489/499
  // type: INFERRED
  // marked bad? no
  // output word of size 10 : index:134 c0nm_b0m_v0m_n247 c0nm_b0m_v0m_n255 c0nm_b0m_v0m_n252 c0nm_b0m_v0m_n251
  // c0nm_b0m_v0m_n250 c0nm_b0m_v0m_n249 c0nm_b0m_v0m_n248 c0nm_b0m_v0m_n246 c0nm_b0m_v0m_n245 c0nm_b0m_v0m_n244
  // group: sel; nodes: [ c0nm_b0m_v0m_n22 c0nm_b0m_v0m_n18 c0nm_b0m_v0m_n20 ]

  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u30 (.A0(c0nm_b0m_v0m_n69), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n70), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n71), .Y(c0nm_b0m_v0m_n244));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u29 (.A0(c0nm_b0m_v0m_n66), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n67), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n68), .Y(c0nm_b0m_v0m_n245));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u28 (.A0(c0nm_b0m_v0m_n63), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n64), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n65), .Y(c0nm_b0m_v0m_n246));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u27 (.A0(c0nm_b0m_v0m_n48), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n49), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n62), .Y(c0nm_b0m_v0m_n247));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u26 (.A0(c0nm_b0m_v0m_n45), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n46), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n47), .Y(c0nm_b0m_v0m_n248));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u25 (.A0(c0nm_b0m_v0m_n42), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n43), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n44), .Y(c0nm_b0m_v0m_n249));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u24 (.A0(c0nm_b0m_v0m_n39), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n40), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n41), .Y(c0nm_b0m_v0m_n250));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u23 (.A0(c0nm_b0m_v0m_n36), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n37), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n38), .Y(c0nm_b0m_v0m_n251));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u22 (.A0(c0nm_b0m_v0m_n33), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n34), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n22), .C1(c0nm_b0m_v0m_n35), .Y(c0nm_b0m_v0m_n252));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u17 (.A0(c0nm_b0m_v0m_n17), .A1(c0nm_b0m_v0m_n18), .B0(c0nm_b0m_v0m_n19), .B1(c0nm_b0m_v0m_n20), .C0(c0nm_b0m_v0m_n21), .C1(c0nm_b0m_v0m_n22), .Y(c0nm_b0m_v0m_n255));
endmodule
module mux31i_oai222_mx27 
(
  c0sm_b0m_v0m_n107, 
  c0sm_b0m_v0m_n129, 
  c0sm_b0m_v0m_n130, 
  c0sm_b0m_v0m_n131, 
  c0sm_b0m_v0m_n138, 
  c0sm_b0m_v0m_n144, 
  c0sm_b0m_v0m_n150, 
  c0sm_b0m_v0m_n156, 
  c0sm_b0m_v0m_n162, 
  c0sm_b0m_v0m_n168, 
  c0sm_b0m_v0m_n17, 
  c0sm_b0m_v0m_n174, 
  c0sm_b0m_v0m_n180, 
  c0sm_b0m_v0m_n186, 
  c0sm_b0m_v0m_n19, 
  c0sm_b0m_v0m_n33, 
  c0sm_b0m_v0m_n34, 
  c0sm_b0m_v0m_n36, 
  c0sm_b0m_v0m_n37, 
  c0sm_b0m_v0m_n39, 
  c0sm_b0m_v0m_n40, 
  c0sm_b0m_v0m_n42, 
  c0sm_b0m_v0m_n43, 
  c0sm_b0m_v0m_n45, 
  c0sm_b0m_v0m_n46, 
  c0sm_b0m_v0m_n48, 
  c0sm_b0m_v0m_n49, 
  c0sm_b0m_v0m_n63, 
  c0sm_b0m_v0m_n64, 
  c0sm_b0m_v0m_n66, 
  c0sm_b0m_v0m_n67, 
  c0sm_b0m_v0m_n69, 
  c0sm_b0m_v0m_n70, 
  c0sm_b0m_v0m_n321,
  c0sm_b0m_v0m_n322,
  c0sm_b0m_v0m_n323,
  c0sm_b0m_v0m_n324,
  c0sm_b0m_v0m_n325,
  c0sm_b0m_v0m_n326,
  c0sm_b0m_v0m_n327,
  c0sm_b0m_v0m_n328,
  c0sm_b0m_v0m_n329,
  c0sm_b0m_v0m_n330
);
  input c0sm_b0m_v0m_n107;
  input c0sm_b0m_v0m_n129;
  input c0sm_b0m_v0m_n130;
  input c0sm_b0m_v0m_n131;
  input c0sm_b0m_v0m_n138;
  input c0sm_b0m_v0m_n144;
  input c0sm_b0m_v0m_n150;
  input c0sm_b0m_v0m_n156;
  input c0sm_b0m_v0m_n162;
  input c0sm_b0m_v0m_n168;
  input c0sm_b0m_v0m_n17;
  input c0sm_b0m_v0m_n174;
  input c0sm_b0m_v0m_n180;
  input c0sm_b0m_v0m_n186;
  input c0sm_b0m_v0m_n19;
  input c0sm_b0m_v0m_n33;
  input c0sm_b0m_v0m_n34;
  input c0sm_b0m_v0m_n36;
  input c0sm_b0m_v0m_n37;
  input c0sm_b0m_v0m_n39;
  input c0sm_b0m_v0m_n40;
  input c0sm_b0m_v0m_n42;
  input c0sm_b0m_v0m_n43;
  input c0sm_b0m_v0m_n45;
  input c0sm_b0m_v0m_n46;
  input c0sm_b0m_v0m_n48;
  input c0sm_b0m_v0m_n49;
  input c0sm_b0m_v0m_n63;
  input c0sm_b0m_v0m_n64;
  input c0sm_b0m_v0m_n66;
  input c0sm_b0m_v0m_n67;
  input c0sm_b0m_v0m_n69;
  input c0sm_b0m_v0m_n70;
  output c0sm_b0m_v0m_n321;
  output c0sm_b0m_v0m_n322;
  output c0sm_b0m_v0m_n323;
  output c0sm_b0m_v0m_n324;
  output c0sm_b0m_v0m_n325;
  output c0sm_b0m_v0m_n326;
  output c0sm_b0m_v0m_n327;
  output c0sm_b0m_v0m_n328;
  output c0sm_b0m_v0m_n329;
  output c0sm_b0m_v0m_n330;

  // moduleNum: x27
  // type: mux31i_oai222
  // conflicting modules: 
  // number of bit inputs: 33
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 500/510
  // type: INFERRED
  // marked bad? no
  // output word of size 10 : index:135 c0sm_b0m_v0m_n321 c0sm_b0m_v0m_n322 c0sm_b0m_v0m_n323 c0sm_b0m_v0m_n324
  // c0sm_b0m_v0m_n325 c0sm_b0m_v0m_n326 c0sm_b0m_v0m_n327 c0sm_b0m_v0m_n328 c0sm_b0m_v0m_n329 c0sm_b0m_v0m_n330
  // group: sel; nodes: [ c0sm_b0m_v0m_n129 c0sm_b0m_v0m_n107 c0sm_b0m_v0m_n130 ]

  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u162 (.A0(c0sm_b0m_v0m_n19), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n17), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n186), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n330));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u155 (.A0(c0sm_b0m_v0m_n70), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n69), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n180), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n329));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u148 (.A0(c0sm_b0m_v0m_n67), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n66), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n174), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n328));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u141 (.A0(c0sm_b0m_v0m_n64), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n63), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n168), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n327));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u134 (.A0(c0sm_b0m_v0m_n49), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n48), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n162), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n326));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u127 (.A0(c0sm_b0m_v0m_n46), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n45), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n156), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n325));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u120 (.A0(c0sm_b0m_v0m_n43), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n42), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n150), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n324));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u113 (.A0(c0sm_b0m_v0m_n40), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n39), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n144), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n323));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u106 (.A0(c0sm_b0m_v0m_n37), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n36), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n138), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n322));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u99 (.A0(c0sm_b0m_v0m_n34), .A1(c0sm_b0m_v0m_n129), .B0(c0sm_b0m_v0m_n33), .B1(c0sm_b0m_v0m_n130), .C0(c0sm_b0m_v0m_n131), .C1(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n321));
endmodule
module mux31i_oai222_mx28 
(
  c0sm_b0m_v0m_n17, 
  c0sm_b0m_v0m_n19, 
  c0sm_b0m_v0m_n33, 
  c0sm_b0m_v0m_n34, 
  c0sm_b0m_v0m_n36, 
  c0sm_b0m_v0m_n37, 
  c0sm_b0m_v0m_n39, 
  c0sm_b0m_v0m_n40, 
  c0sm_b0m_v0m_n42, 
  c0sm_b0m_v0m_n43, 
  c0sm_b0m_v0m_n45, 
  c0sm_b0m_v0m_n46, 
  c0sm_b0m_v0m_n48, 
  c0sm_b0m_v0m_n49, 
  c0sm_b0m_v0m_n63, 
  c0sm_b0m_v0m_n64, 
  c0sm_b0m_v0m_n66, 
  c0sm_b0m_v0m_n67, 
  c0sm_b0m_v0m_n69, 
  c0sm_b0m_v0m_n70, 
  c0sm_b0m_v0m_n76, 
  c0sm_b0m_v0m_n81, 
  c0sm_b0m_v0m_n82, 
  c0sm_b0m_v0m_n83, 
  c0sm_b0m_v0m_n84, 
  c0sm_b0m_v0m_n85, 
  c0sm_b0m_v0m_n86, 
  c0sm_b0m_v0m_n87, 
  c0sm_b0m_v0m_n88, 
  c0sm_b0m_v0m_n89, 
  c0sm_b0m_v0m_n90, 
  c0sm_b0m_v0m_n91, 
  c0sm_b0m_v0m_n92, 
  c0sm_b0m_v0m_n297,
  c0sm_b0m_v0m_n298,
  c0sm_b0m_v0m_n299,
  c0sm_b0m_v0m_n300,
  c0sm_b0m_v0m_n301,
  c0sm_b0m_v0m_n302,
  c0sm_b0m_v0m_n303,
  c0sm_b0m_v0m_n304,
  c0sm_b0m_v0m_n305,
  c0sm_b0m_v0m_n306
);
  input c0sm_b0m_v0m_n17;
  input c0sm_b0m_v0m_n19;
  input c0sm_b0m_v0m_n33;
  input c0sm_b0m_v0m_n34;
  input c0sm_b0m_v0m_n36;
  input c0sm_b0m_v0m_n37;
  input c0sm_b0m_v0m_n39;
  input c0sm_b0m_v0m_n40;
  input c0sm_b0m_v0m_n42;
  input c0sm_b0m_v0m_n43;
  input c0sm_b0m_v0m_n45;
  input c0sm_b0m_v0m_n46;
  input c0sm_b0m_v0m_n48;
  input c0sm_b0m_v0m_n49;
  input c0sm_b0m_v0m_n63;
  input c0sm_b0m_v0m_n64;
  input c0sm_b0m_v0m_n66;
  input c0sm_b0m_v0m_n67;
  input c0sm_b0m_v0m_n69;
  input c0sm_b0m_v0m_n70;
  input c0sm_b0m_v0m_n76;
  input c0sm_b0m_v0m_n81;
  input c0sm_b0m_v0m_n82;
  input c0sm_b0m_v0m_n83;
  input c0sm_b0m_v0m_n84;
  input c0sm_b0m_v0m_n85;
  input c0sm_b0m_v0m_n86;
  input c0sm_b0m_v0m_n87;
  input c0sm_b0m_v0m_n88;
  input c0sm_b0m_v0m_n89;
  input c0sm_b0m_v0m_n90;
  input c0sm_b0m_v0m_n91;
  input c0sm_b0m_v0m_n92;
  output c0sm_b0m_v0m_n297;
  output c0sm_b0m_v0m_n298;
  output c0sm_b0m_v0m_n299;
  output c0sm_b0m_v0m_n300;
  output c0sm_b0m_v0m_n301;
  output c0sm_b0m_v0m_n302;
  output c0sm_b0m_v0m_n303;
  output c0sm_b0m_v0m_n304;
  output c0sm_b0m_v0m_n305;
  output c0sm_b0m_v0m_n306;

  // moduleNum: x28
  // type: mux31i_oai222
  // conflicting modules: 
  // number of bit inputs: 33
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 522/532
  // type: INFERRED
  // marked bad? no
  // output word of size 10 : index:137 c0sm_b0m_v0m_n301 c0sm_b0m_v0m_n300 c0sm_b0m_v0m_n299 c0sm_b0m_v0m_n298
  // c0sm_b0m_v0m_n297 c0sm_b0m_v0m_n302 c0sm_b0m_v0m_n305 c0sm_b0m_v0m_n306 c0sm_b0m_v0m_n304 c0sm_b0m_v0m_n303
  // group: sel; nodes: [ c0sm_b0m_v0m_n81 c0sm_b0m_v0m_n76 c0sm_b0m_v0m_n82 ]

  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u58 (.A0(c0sm_b0m_v0m_n19), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n17), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n92), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n306));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u56 (.A0(c0sm_b0m_v0m_n70), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n69), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n91), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n305));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u54 (.A0(c0sm_b0m_v0m_n67), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n66), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n90), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n304));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u52 (.A0(c0sm_b0m_v0m_n64), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n63), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n89), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n303));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u50 (.A0(c0sm_b0m_v0m_n49), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n48), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n88), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n302));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u48 (.A0(c0sm_b0m_v0m_n46), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n45), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n87), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n301));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u46 (.A0(c0sm_b0m_v0m_n43), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n42), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n86), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n300));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u44 (.A0(c0sm_b0m_v0m_n40), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n39), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n85), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n299));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u42 (.A0(c0sm_b0m_v0m_n37), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n36), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n84), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n298));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u40 (.A0(c0sm_b0m_v0m_n34), .A1(c0sm_b0m_v0m_n81), .B0(c0sm_b0m_v0m_n33), .B1(c0sm_b0m_v0m_n82), .C0(c0sm_b0m_v0m_n83), .C1(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n297));
endmodule
module mux31i_oai222_mx29 
(
  c0sm_b0m_v0m_n17, 
  c0sm_b0m_v0m_n18, 
  c0sm_b0m_v0m_n19, 
  c0sm_b0m_v0m_n20, 
  c0sm_b0m_v0m_n21, 
  c0sm_b0m_v0m_n22, 
  c0sm_b0m_v0m_n33, 
  c0sm_b0m_v0m_n34, 
  c0sm_b0m_v0m_n35, 
  c0sm_b0m_v0m_n36, 
  c0sm_b0m_v0m_n37, 
  c0sm_b0m_v0m_n38, 
  c0sm_b0m_v0m_n39, 
  c0sm_b0m_v0m_n40, 
  c0sm_b0m_v0m_n41, 
  c0sm_b0m_v0m_n42, 
  c0sm_b0m_v0m_n43, 
  c0sm_b0m_v0m_n44, 
  c0sm_b0m_v0m_n45, 
  c0sm_b0m_v0m_n46, 
  c0sm_b0m_v0m_n47, 
  c0sm_b0m_v0m_n48, 
  c0sm_b0m_v0m_n49, 
  c0sm_b0m_v0m_n62, 
  c0sm_b0m_v0m_n63, 
  c0sm_b0m_v0m_n64, 
  c0sm_b0m_v0m_n65, 
  c0sm_b0m_v0m_n66, 
  c0sm_b0m_v0m_n67, 
  c0sm_b0m_v0m_n68, 
  c0sm_b0m_v0m_n69, 
  c0sm_b0m_v0m_n70, 
  c0sm_b0m_v0m_n71, 
  c0sm_b0m_v0m_n283,
  c0sm_b0m_v0m_n286,
  c0sm_b0m_v0m_n287,
  c0sm_b0m_v0m_n288,
  c0sm_b0m_v0m_n289,
  c0sm_b0m_v0m_n290,
  c0sm_b0m_v0m_n291,
  c0sm_b0m_v0m_n292,
  c0sm_b0m_v0m_n293,
  c0sm_b0m_v0m_n294
);
  input c0sm_b0m_v0m_n17;
  input c0sm_b0m_v0m_n18;
  input c0sm_b0m_v0m_n19;
  input c0sm_b0m_v0m_n20;
  input c0sm_b0m_v0m_n21;
  input c0sm_b0m_v0m_n22;
  input c0sm_b0m_v0m_n33;
  input c0sm_b0m_v0m_n34;
  input c0sm_b0m_v0m_n35;
  input c0sm_b0m_v0m_n36;
  input c0sm_b0m_v0m_n37;
  input c0sm_b0m_v0m_n38;
  input c0sm_b0m_v0m_n39;
  input c0sm_b0m_v0m_n40;
  input c0sm_b0m_v0m_n41;
  input c0sm_b0m_v0m_n42;
  input c0sm_b0m_v0m_n43;
  input c0sm_b0m_v0m_n44;
  input c0sm_b0m_v0m_n45;
  input c0sm_b0m_v0m_n46;
  input c0sm_b0m_v0m_n47;
  input c0sm_b0m_v0m_n48;
  input c0sm_b0m_v0m_n49;
  input c0sm_b0m_v0m_n62;
  input c0sm_b0m_v0m_n63;
  input c0sm_b0m_v0m_n64;
  input c0sm_b0m_v0m_n65;
  input c0sm_b0m_v0m_n66;
  input c0sm_b0m_v0m_n67;
  input c0sm_b0m_v0m_n68;
  input c0sm_b0m_v0m_n69;
  input c0sm_b0m_v0m_n70;
  input c0sm_b0m_v0m_n71;
  output c0sm_b0m_v0m_n283;
  output c0sm_b0m_v0m_n286;
  output c0sm_b0m_v0m_n287;
  output c0sm_b0m_v0m_n288;
  output c0sm_b0m_v0m_n289;
  output c0sm_b0m_v0m_n290;
  output c0sm_b0m_v0m_n291;
  output c0sm_b0m_v0m_n292;
  output c0sm_b0m_v0m_n293;
  output c0sm_b0m_v0m_n294;

  // moduleNum: x29
  // type: mux31i_oai222
  // conflicting modules: 
  // number of bit inputs: 33
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 533/543
  // type: INFERRED
  // marked bad? no
  // output word of size 10 : index:138 c0sm_b0m_v0m_n288 c0sm_b0m_v0m_n294 c0sm_b0m_v0m_n293 c0sm_b0m_v0m_n292
  // c0sm_b0m_v0m_n291 c0sm_b0m_v0m_n290 c0sm_b0m_v0m_n289 c0sm_b0m_v0m_n287 c0sm_b0m_v0m_n286 c0sm_b0m_v0m_n283
  // group: sel; nodes: [ c0sm_b0m_v0m_n22 c0sm_b0m_v0m_n18 c0sm_b0m_v0m_n20 ]

  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u30 (.A0(c0sm_b0m_v0m_n69), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n70), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n71), .Y(c0sm_b0m_v0m_n294));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u29 (.A0(c0sm_b0m_v0m_n66), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n67), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n68), .Y(c0sm_b0m_v0m_n293));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u28 (.A0(c0sm_b0m_v0m_n63), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n64), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n65), .Y(c0sm_b0m_v0m_n292));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u27 (.A0(c0sm_b0m_v0m_n48), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n49), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n62), .Y(c0sm_b0m_v0m_n291));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u26 (.A0(c0sm_b0m_v0m_n45), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n46), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n47), .Y(c0sm_b0m_v0m_n290));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u25 (.A0(c0sm_b0m_v0m_n42), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n43), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n44), .Y(c0sm_b0m_v0m_n289));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u24 (.A0(c0sm_b0m_v0m_n39), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n40), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n41), .Y(c0sm_b0m_v0m_n288));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u23 (.A0(c0sm_b0m_v0m_n36), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n37), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n38), .Y(c0sm_b0m_v0m_n287));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u22 (.A0(c0sm_b0m_v0m_n33), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n34), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n22), .C1(c0sm_b0m_v0m_n35), .Y(c0sm_b0m_v0m_n286));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u17 (.A0(c0sm_b0m_v0m_n17), .A1(c0sm_b0m_v0m_n18), .B0(c0sm_b0m_v0m_n19), .B1(c0sm_b0m_v0m_n20), .C0(c0sm_b0m_v0m_n21), .C1(c0sm_b0m_v0m_n22), .Y(c0sm_b0m_v0m_n283));
endmodule
module mux21i_aoi221_mx30 
(
  c0nm_r0m_n10, 
  c0nm_r0m_n8, 
  c0nm_r0m_n9, 
  c0sm_r0m_n10, 
  c0sm_r0m_n8, 
  c0sm_r0m_n9, 
  currx_0_, 
  currx_1_, 
  c0nm_r0m_n7,
  c0sm_r0m_n7
);
  input c0nm_r0m_n10;
  input c0nm_r0m_n8;
  input c0nm_r0m_n9;
  input c0sm_r0m_n10;
  input c0sm_r0m_n8;
  input c0sm_r0m_n9;
  input currx_0_;
  input currx_1_;
  output c0nm_r0m_n7;
  output c0sm_r0m_n7;

  // moduleNum: x30
  // type: mux21i_aoi221
  // conflicting modules: 
  // number of bit inputs: 8
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 544/544
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:139 c0sm_r0m_n7 c0nm_r0m_n7 
  // group: sel; nodes: [ currx[1] currx[0] ]

  AOI221_X0P5M_A12TR c0nm_r0m_u9 (.A0(currx_1_), .A1(c0nm_r0m_n8), .B0(currx_0_), .B1(c0nm_r0m_n9), .C0(c0nm_r0m_n10), .Y(c0nm_r0m_n7));
  AOI221_X0P5M_A12TR c0sm_r0m_u9 (.A0(currx_1_), .A1(c0sm_r0m_n8), .B0(currx_0_), .B1(c0sm_r0m_n9), .C0(c0sm_r0m_n10), .Y(c0sm_r0m_n7));
endmodule
module mux21i_aoi221_mx31 
(
  c0sm_b0m_v0m_n100, 
  c0sm_b0m_v0m_n25, 
  c0sm_b0m_v0m_n27, 
  c0sm_b0m_v0m_n31, 
  c0sm_b0m_v0m_n32, 
  c0sm_b0m_v0m_n99, 
  reset, 
  c0sm_b0m_v0m_n101,
  c0sm_b0m_v0m_n97
);
  input c0sm_b0m_v0m_n100;
  input c0sm_b0m_v0m_n25;
  input c0sm_b0m_v0m_n27;
  input c0sm_b0m_v0m_n31;
  input c0sm_b0m_v0m_n32;
  input c0sm_b0m_v0m_n99;
  input reset;
  output c0sm_b0m_v0m_n101;
  output c0sm_b0m_v0m_n97;

  // moduleNum: x31
  // type: mux21i_aoi221
  // conflicting modules: 
  // number of bit inputs: 7
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 624/626
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:-1 c0sm_b0m_v0m_n101 c0sm_b0m_v0m_n97 
  // group: sel; nodes: [ reset c0sm_b0m_v0m_n100 ]

  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u68 (.A0(c0sm_b0m_v0m_n99), .A1(c0sm_b0m_v0m_n31), .B0(c0sm_b0m_v0m_n100), .B1(c0sm_b0m_v0m_n32), .C0(reset), .Y(c0sm_b0m_v0m_n101));
  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u66 (.A0(c0sm_b0m_v0m_n99), .A1(c0sm_b0m_v0m_n25), .B0(c0sm_b0m_v0m_n100), .B1(c0sm_b0m_v0m_n27), .C0(reset), .Y(c0sm_b0m_v0m_n97));
endmodule
module mux21i_aoi221_mx32 
(
  c0nm_b0m_v0m_n100, 
  c0nm_b0m_v0m_n25, 
  c0nm_b0m_v0m_n27, 
  c0nm_b0m_v0m_n31, 
  c0nm_b0m_v0m_n32, 
  c0nm_b0m_v0m_n99, 
  reset, 
  c0nm_b0m_v0m_n101,
  c0nm_b0m_v0m_n97
);
  input c0nm_b0m_v0m_n100;
  input c0nm_b0m_v0m_n25;
  input c0nm_b0m_v0m_n27;
  input c0nm_b0m_v0m_n31;
  input c0nm_b0m_v0m_n32;
  input c0nm_b0m_v0m_n99;
  input reset;
  output c0nm_b0m_v0m_n101;
  output c0nm_b0m_v0m_n97;

  // moduleNum: x32
  // type: mux21i_aoi221
  // conflicting modules: 
  // number of bit inputs: 7
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 749/751
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:-1 c0nm_b0m_v0m_n101 c0nm_b0m_v0m_n97 
  // group: sel; nodes: [ c0nm_b0m_v0m_n99 c0nm_b0m_v0m_n100 ]

  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u68 (.A0(c0nm_b0m_v0m_n99), .A1(c0nm_b0m_v0m_n31), .B0(c0nm_b0m_v0m_n100), .B1(c0nm_b0m_v0m_n32), .C0(reset), .Y(c0nm_b0m_v0m_n101));
  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u66 (.A0(c0nm_b0m_v0m_n99), .A1(c0nm_b0m_v0m_n25), .B0(c0nm_b0m_v0m_n100), .B1(c0nm_b0m_v0m_n27), .C0(reset), .Y(c0nm_b0m_v0m_n97));
endmodule
module mux21i_aoi221_mx33 
(
  c0sm_b0m_v0m_buffers0_0_, 
  c0sm_b0m_v0m_buffers0_1_, 
  c0sm_b0m_v0m_n113, 
  c0sm_b0m_v0m_n114, 
  c0sm_b0m_v0m_n115, 
  c0sm_b0m_v0m_n125, 
  debitout_1, 
  c0sm_b0m_v0m_n112,
  c0sm_b0m_v0m_n124
);
  input c0sm_b0m_v0m_buffers0_0_;
  input c0sm_b0m_v0m_buffers0_1_;
  input c0sm_b0m_v0m_n113;
  input c0sm_b0m_v0m_n114;
  input c0sm_b0m_v0m_n115;
  input c0sm_b0m_v0m_n125;
  input debitout_1;
  output c0sm_b0m_v0m_n112;
  output c0sm_b0m_v0m_n124;

  // moduleNum: x33
  // type: mux21i_aoi221
  // conflicting modules: 
  // number of bit inputs: 7
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 846/848
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:-1 c0sm_b0m_v0m_n112 c0sm_b0m_v0m_n124 
  // group: sel; nodes: [ c0sm_b0m_v0m_n115 c0sm_b0m_v0m_n113 ]

  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u94 (.A0(c0sm_b0m_v0m_n113), .A1(c0sm_b0m_v0m_n125), .B0(c0sm_b0m_v0m_buffers0_1_), .B1(c0sm_b0m_v0m_n115), .C0(debitout_1), .Y(c0sm_b0m_v0m_n124));
  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u87 (.A0(c0sm_b0m_v0m_n113), .A1(c0sm_b0m_v0m_n114), .B0(c0sm_b0m_v0m_buffers0_0_), .B1(c0sm_b0m_v0m_n115), .C0(debitout_1), .Y(c0sm_b0m_v0m_n112));
endmodule
module mux21_oa221_mx34 
(
  c0nm_b0m_v0m_n138, 
  c0nm_b0m_v0m_n150, 
  c0nm_b0m_v0m_n156, 
  c0nm_b0m_v0m_n187, 
  c0nm_b0m_v0m_n268, 
  c0nm_b0m_v0m_n269, 
  c0nm_b0m_v0m_n271, 
  c0nm_b0m_v0m_n38, 
  c0nm_b0m_v0m_n44, 
  c0nm_b0m_v0m_n47, 
  c0nm_b0m_v0m_n73, 
  c0nm_r0m_n14,
  c0nm_r0m_n8,
  c0nm_r0m_n9
);
  input c0nm_b0m_v0m_n138;
  input c0nm_b0m_v0m_n150;
  input c0nm_b0m_v0m_n156;
  input c0nm_b0m_v0m_n187;
  input c0nm_b0m_v0m_n268;
  input c0nm_b0m_v0m_n269;
  input c0nm_b0m_v0m_n271;
  input c0nm_b0m_v0m_n38;
  input c0nm_b0m_v0m_n44;
  input c0nm_b0m_v0m_n47;
  input c0nm_b0m_v0m_n73;
  output c0nm_r0m_n14;
  output c0nm_r0m_n8;
  output c0nm_r0m_n9;
  wire c0nm_headflit_3_;
  wire c0nm_headflit_5_;
  wire c0nm_headflit_6_;

  // moduleNum: x34
  // type: mux21_oa221
  // conflicting modules: 
  // number of bit inputs: 11
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 6
  // number of non-inferred gates: 0
  // ILP vars: 897/901
  // type: INFERRED
  // marked bad? no
  // output word of size 3 : index:243 c0nm_r0m_n14 c0nm_r0m_n8 c0nm_r0m_n9 
  // group: sel; nodes: [ c0nm_b0m_v0m_n187 c0nm_b0m_v0m_n73 ]

  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u240 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n138), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n38), .C0(c0nm_b0m_v0m_n271), .Y(c0nm_headflit_3_));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u230 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n150), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n44), .C0(c0nm_b0m_v0m_n269), .Y(c0nm_headflit_5_));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u225 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n156), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n47), .C0(c0nm_b0m_v0m_n268), .Y(c0nm_headflit_6_));
  INV_X0P5B_A12TR c0nm_r0m_u19 (.A(c0nm_headflit_5_), .Y(c0nm_r0m_n9));
  INV_X0P5B_A12TR c0nm_r0m_u17 (.A(c0nm_headflit_6_), .Y(c0nm_r0m_n8));
  INV_X0P5B_A12TR c0nm_r0m_u13 (.A(c0nm_headflit_3_), .Y(c0nm_r0m_n14));
endmodule
module mux21_oa221_mx35 
(
  c0nm_b0m_v0m_n110, 
  c0nm_b0m_v0m_n111, 
  c0nm_b0m_v0m_n131, 
  c0nm_b0m_v0m_n133, 
  c0nm_b0m_v0m_n138, 
  c0nm_b0m_v0m_n140, 
  c0nm_b0m_v0m_n144, 
  c0nm_b0m_v0m_n146, 
  c0nm_b0m_v0m_n150, 
  c0nm_b0m_v0m_n152, 
  c0nm_b0m_v0m_n156, 
  c0nm_b0m_v0m_n158, 
  c0nm_b0m_v0m_n162, 
  c0nm_b0m_v0m_n164, 
  c0nm_b0m_v0m_n168, 
  c0nm_b0m_v0m_n170, 
  c0nm_b0m_v0m_n174, 
  c0nm_b0m_v0m_n176, 
  c0nm_b0m_v0m_n180, 
  c0nm_b0m_v0m_n182, 
  c0nm_b0m_v0m_n186, 
  c0nm_b0m_v0m_n189, 
  c0nm_b0m_v0m_n21, 
  c0nm_b0m_v0m_n35, 
  c0nm_b0m_v0m_n38, 
  c0nm_b0m_v0m_n41, 
  c0nm_b0m_v0m_n44, 
  c0nm_b0m_v0m_n47, 
  c0nm_b0m_v0m_n62, 
  c0nm_b0m_v0m_n65, 
  c0nm_b0m_v0m_n68, 
  c0nm_b0m_v0m_n71, 
  c0nm_b0m_v0m_n17,
  c0nm_b0m_v0m_n33,
  c0nm_b0m_v0m_n36,
  c0nm_b0m_v0m_n39,
  c0nm_b0m_v0m_n42,
  c0nm_b0m_v0m_n45,
  c0nm_b0m_v0m_n48,
  c0nm_b0m_v0m_n63,
  c0nm_b0m_v0m_n66,
  c0nm_b0m_v0m_n69
);
  input c0nm_b0m_v0m_n110;
  input c0nm_b0m_v0m_n111;
  input c0nm_b0m_v0m_n131;
  input c0nm_b0m_v0m_n133;
  input c0nm_b0m_v0m_n138;
  input c0nm_b0m_v0m_n140;
  input c0nm_b0m_v0m_n144;
  input c0nm_b0m_v0m_n146;
  input c0nm_b0m_v0m_n150;
  input c0nm_b0m_v0m_n152;
  input c0nm_b0m_v0m_n156;
  input c0nm_b0m_v0m_n158;
  input c0nm_b0m_v0m_n162;
  input c0nm_b0m_v0m_n164;
  input c0nm_b0m_v0m_n168;
  input c0nm_b0m_v0m_n170;
  input c0nm_b0m_v0m_n174;
  input c0nm_b0m_v0m_n176;
  input c0nm_b0m_v0m_n180;
  input c0nm_b0m_v0m_n182;
  input c0nm_b0m_v0m_n186;
  input c0nm_b0m_v0m_n189;
  input c0nm_b0m_v0m_n21;
  input c0nm_b0m_v0m_n35;
  input c0nm_b0m_v0m_n38;
  input c0nm_b0m_v0m_n41;
  input c0nm_b0m_v0m_n44;
  input c0nm_b0m_v0m_n47;
  input c0nm_b0m_v0m_n62;
  input c0nm_b0m_v0m_n65;
  input c0nm_b0m_v0m_n68;
  input c0nm_b0m_v0m_n71;
  output c0nm_b0m_v0m_n17;
  output c0nm_b0m_v0m_n33;
  output c0nm_b0m_v0m_n36;
  output c0nm_b0m_v0m_n39;
  output c0nm_b0m_v0m_n42;
  output c0nm_b0m_v0m_n45;
  output c0nm_b0m_v0m_n48;
  output c0nm_b0m_v0m_n63;
  output c0nm_b0m_v0m_n66;
  output c0nm_b0m_v0m_n69;
  wire c0nm_b0m_v0m_n132;
  wire c0nm_b0m_v0m_n139;
  wire c0nm_b0m_v0m_n145;
  wire c0nm_b0m_v0m_n151;
  wire c0nm_b0m_v0m_n157;
  wire c0nm_b0m_v0m_n163;
  wire c0nm_b0m_v0m_n169;
  wire c0nm_b0m_v0m_n175;
  wire c0nm_b0m_v0m_n181;
  wire c0nm_b0m_v0m_n188;

  // moduleNum: x35
  // type: mux21_oa221
  // conflicting modules: 
  // number of bit inputs: 32
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 20
  // number of non-inferred gates: 0
  // ILP vars: 911/921
  // type: INFERRED
  // marked bad? no
  // output word of size 10 : index:162 c0nm_b0m_v0m_n33 c0nm_b0m_v0m_n36 c0nm_b0m_v0m_n69 c0nm_b0m_v0m_n66 c0nm_b0m_v0m_n39
  // c0nm_b0m_v0m_n42 c0nm_b0m_v0m_n63 c0nm_b0m_v0m_n48 c0nm_b0m_v0m_n45 c0nm_b0m_v0m_n17
  // group: sel; nodes: [ c0nm_b0m_v0m_n111 c0nm_b0m_v0m_n110 ]

  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u169 (.A0(c0nm_b0m_v0m_n21), .A1(c0nm_b0m_v0m_n111), .B0(c0nm_b0m_v0m_n186), .B1(c0nm_b0m_v0m_n110), .C0(c0nm_b0m_v0m_n189), .Y(c0nm_b0m_v0m_n188));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u168 (.A(c0nm_b0m_v0m_n188), .Y(c0nm_b0m_v0m_n17));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u157 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n71), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n180), .C0(c0nm_b0m_v0m_n182), .Y(c0nm_b0m_v0m_n181));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u156 (.A(c0nm_b0m_v0m_n181), .Y(c0nm_b0m_v0m_n69));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u150 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n68), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n174), .C0(c0nm_b0m_v0m_n176), .Y(c0nm_b0m_v0m_n175));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u149 (.A(c0nm_b0m_v0m_n175), .Y(c0nm_b0m_v0m_n66));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u143 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n65), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n168), .C0(c0nm_b0m_v0m_n170), .Y(c0nm_b0m_v0m_n169));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u142 (.A(c0nm_b0m_v0m_n169), .Y(c0nm_b0m_v0m_n63));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u136 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n62), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n162), .C0(c0nm_b0m_v0m_n164), .Y(c0nm_b0m_v0m_n163));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u135 (.A(c0nm_b0m_v0m_n163), .Y(c0nm_b0m_v0m_n48));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u129 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n47), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n156), .C0(c0nm_b0m_v0m_n158), .Y(c0nm_b0m_v0m_n157));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u128 (.A(c0nm_b0m_v0m_n157), .Y(c0nm_b0m_v0m_n45));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u122 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n44), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n150), .C0(c0nm_b0m_v0m_n152), .Y(c0nm_b0m_v0m_n151));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u121 (.A(c0nm_b0m_v0m_n151), .Y(c0nm_b0m_v0m_n42));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u115 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n41), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n144), .C0(c0nm_b0m_v0m_n146), .Y(c0nm_b0m_v0m_n145));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u114 (.A(c0nm_b0m_v0m_n145), .Y(c0nm_b0m_v0m_n39));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u108 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n38), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n138), .C0(c0nm_b0m_v0m_n140), .Y(c0nm_b0m_v0m_n139));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u107 (.A(c0nm_b0m_v0m_n139), .Y(c0nm_b0m_v0m_n36));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u101 (.A0(c0nm_b0m_v0m_n111), .A1(c0nm_b0m_v0m_n35), .B0(c0nm_b0m_v0m_n110), .B1(c0nm_b0m_v0m_n131), .C0(c0nm_b0m_v0m_n133), .Y(c0nm_b0m_v0m_n132));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u100 (.A(c0nm_b0m_v0m_n132), .Y(c0nm_b0m_v0m_n33));
endmodule
module mux21_oa221_mx36 
(
  c0sm_b0m_v0m_n138, 
  c0sm_b0m_v0m_n150, 
  c0sm_b0m_v0m_n156, 
  c0sm_b0m_v0m_n187, 
  c0sm_b0m_v0m_n268, 
  c0sm_b0m_v0m_n269, 
  c0sm_b0m_v0m_n271, 
  c0sm_b0m_v0m_n38, 
  c0sm_b0m_v0m_n44, 
  c0sm_b0m_v0m_n47, 
  c0sm_b0m_v0m_n73, 
  c0sm_r0m_n14,
  c0sm_r0m_n8,
  c0sm_r0m_n9
);
  input c0sm_b0m_v0m_n138;
  input c0sm_b0m_v0m_n150;
  input c0sm_b0m_v0m_n156;
  input c0sm_b0m_v0m_n187;
  input c0sm_b0m_v0m_n268;
  input c0sm_b0m_v0m_n269;
  input c0sm_b0m_v0m_n271;
  input c0sm_b0m_v0m_n38;
  input c0sm_b0m_v0m_n44;
  input c0sm_b0m_v0m_n47;
  input c0sm_b0m_v0m_n73;
  output c0sm_r0m_n14;
  output c0sm_r0m_n8;
  output c0sm_r0m_n9;
  wire c0sm_headflit_3_;
  wire c0sm_headflit_5_;
  wire c0sm_headflit_6_;

  // moduleNum: x36
  // type: mux21_oa221
  // conflicting modules: 
  // number of bit inputs: 11
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 6
  // number of non-inferred gates: 0
  // ILP vars: 922/926
  // type: INFERRED
  // marked bad? no
  // output word of size 3 : index:244 c0sm_r0m_n14 c0sm_r0m_n9 c0sm_r0m_n8 
  // group: sel; nodes: [ c0sm_b0m_v0m_n187 c0sm_b0m_v0m_n73 ]

  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u240 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n138), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n38), .C0(c0sm_b0m_v0m_n271), .Y(c0sm_headflit_3_));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u230 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n150), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n44), .C0(c0sm_b0m_v0m_n269), .Y(c0sm_headflit_5_));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u225 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n156), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n47), .C0(c0sm_b0m_v0m_n268), .Y(c0sm_headflit_6_));
  INV_X0P5B_A12TR c0sm_r0m_u19 (.A(c0sm_headflit_5_), .Y(c0sm_r0m_n9));
  INV_X0P5B_A12TR c0sm_r0m_u17 (.A(c0sm_headflit_6_), .Y(c0sm_r0m_n8));
  INV_X0P5B_A12TR c0sm_r0m_u13 (.A(c0sm_headflit_3_), .Y(c0sm_r0m_n14));
endmodule
module mux21_oa221_mx37 
(
  c0sm_b0m_v0m_n110, 
  c0sm_b0m_v0m_n111, 
  c0sm_b0m_v0m_n131, 
  c0sm_b0m_v0m_n133, 
  c0sm_b0m_v0m_n138, 
  c0sm_b0m_v0m_n140, 
  c0sm_b0m_v0m_n144, 
  c0sm_b0m_v0m_n146, 
  c0sm_b0m_v0m_n150, 
  c0sm_b0m_v0m_n152, 
  c0sm_b0m_v0m_n156, 
  c0sm_b0m_v0m_n158, 
  c0sm_b0m_v0m_n162, 
  c0sm_b0m_v0m_n164, 
  c0sm_b0m_v0m_n168, 
  c0sm_b0m_v0m_n170, 
  c0sm_b0m_v0m_n174, 
  c0sm_b0m_v0m_n176, 
  c0sm_b0m_v0m_n180, 
  c0sm_b0m_v0m_n182, 
  c0sm_b0m_v0m_n186, 
  c0sm_b0m_v0m_n189, 
  c0sm_b0m_v0m_n21, 
  c0sm_b0m_v0m_n35, 
  c0sm_b0m_v0m_n38, 
  c0sm_b0m_v0m_n41, 
  c0sm_b0m_v0m_n44, 
  c0sm_b0m_v0m_n47, 
  c0sm_b0m_v0m_n62, 
  c0sm_b0m_v0m_n65, 
  c0sm_b0m_v0m_n68, 
  c0sm_b0m_v0m_n71, 
  c0sm_b0m_v0m_n17,
  c0sm_b0m_v0m_n33,
  c0sm_b0m_v0m_n36,
  c0sm_b0m_v0m_n39,
  c0sm_b0m_v0m_n42,
  c0sm_b0m_v0m_n45,
  c0sm_b0m_v0m_n48,
  c0sm_b0m_v0m_n63,
  c0sm_b0m_v0m_n66,
  c0sm_b0m_v0m_n69
);
  input c0sm_b0m_v0m_n110;
  input c0sm_b0m_v0m_n111;
  input c0sm_b0m_v0m_n131;
  input c0sm_b0m_v0m_n133;
  input c0sm_b0m_v0m_n138;
  input c0sm_b0m_v0m_n140;
  input c0sm_b0m_v0m_n144;
  input c0sm_b0m_v0m_n146;
  input c0sm_b0m_v0m_n150;
  input c0sm_b0m_v0m_n152;
  input c0sm_b0m_v0m_n156;
  input c0sm_b0m_v0m_n158;
  input c0sm_b0m_v0m_n162;
  input c0sm_b0m_v0m_n164;
  input c0sm_b0m_v0m_n168;
  input c0sm_b0m_v0m_n170;
  input c0sm_b0m_v0m_n174;
  input c0sm_b0m_v0m_n176;
  input c0sm_b0m_v0m_n180;
  input c0sm_b0m_v0m_n182;
  input c0sm_b0m_v0m_n186;
  input c0sm_b0m_v0m_n189;
  input c0sm_b0m_v0m_n21;
  input c0sm_b0m_v0m_n35;
  input c0sm_b0m_v0m_n38;
  input c0sm_b0m_v0m_n41;
  input c0sm_b0m_v0m_n44;
  input c0sm_b0m_v0m_n47;
  input c0sm_b0m_v0m_n62;
  input c0sm_b0m_v0m_n65;
  input c0sm_b0m_v0m_n68;
  input c0sm_b0m_v0m_n71;
  output c0sm_b0m_v0m_n17;
  output c0sm_b0m_v0m_n33;
  output c0sm_b0m_v0m_n36;
  output c0sm_b0m_v0m_n39;
  output c0sm_b0m_v0m_n42;
  output c0sm_b0m_v0m_n45;
  output c0sm_b0m_v0m_n48;
  output c0sm_b0m_v0m_n63;
  output c0sm_b0m_v0m_n66;
  output c0sm_b0m_v0m_n69;
  wire c0sm_b0m_v0m_n132;
  wire c0sm_b0m_v0m_n139;
  wire c0sm_b0m_v0m_n145;
  wire c0sm_b0m_v0m_n151;
  wire c0sm_b0m_v0m_n157;
  wire c0sm_b0m_v0m_n163;
  wire c0sm_b0m_v0m_n169;
  wire c0sm_b0m_v0m_n175;
  wire c0sm_b0m_v0m_n181;
  wire c0sm_b0m_v0m_n188;

  // moduleNum: x37
  // type: mux21_oa221
  // conflicting modules: 
  // number of bit inputs: 32
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 20
  // number of non-inferred gates: 0
  // ILP vars: 936/946
  // type: INFERRED
  // marked bad? no
  // output word of size 10 : index:167 c0sm_b0m_v0m_n33 c0sm_b0m_v0m_n48 c0sm_b0m_v0m_n17 c0sm_b0m_v0m_n45 c0sm_b0m_v0m_n42
  // c0sm_b0m_v0m_n63 c0sm_b0m_v0m_n66 c0sm_b0m_v0m_n39 c0sm_b0m_v0m_n69 c0sm_b0m_v0m_n36
  // group: sel; nodes: [ c0sm_b0m_v0m_n111 c0sm_b0m_v0m_n110 ]

  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u169 (.A0(c0sm_b0m_v0m_n21), .A1(c0sm_b0m_v0m_n111), .B0(c0sm_b0m_v0m_n186), .B1(c0sm_b0m_v0m_n110), .C0(c0sm_b0m_v0m_n189), .Y(c0sm_b0m_v0m_n188));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u168 (.A(c0sm_b0m_v0m_n188), .Y(c0sm_b0m_v0m_n17));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u157 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n71), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n180), .C0(c0sm_b0m_v0m_n182), .Y(c0sm_b0m_v0m_n181));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u156 (.A(c0sm_b0m_v0m_n181), .Y(c0sm_b0m_v0m_n69));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u150 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n68), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n174), .C0(c0sm_b0m_v0m_n176), .Y(c0sm_b0m_v0m_n175));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u149 (.A(c0sm_b0m_v0m_n175), .Y(c0sm_b0m_v0m_n66));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u143 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n65), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n168), .C0(c0sm_b0m_v0m_n170), .Y(c0sm_b0m_v0m_n169));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u142 (.A(c0sm_b0m_v0m_n169), .Y(c0sm_b0m_v0m_n63));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u136 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n62), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n162), .C0(c0sm_b0m_v0m_n164), .Y(c0sm_b0m_v0m_n163));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u135 (.A(c0sm_b0m_v0m_n163), .Y(c0sm_b0m_v0m_n48));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u129 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n47), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n156), .C0(c0sm_b0m_v0m_n158), .Y(c0sm_b0m_v0m_n157));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u128 (.A(c0sm_b0m_v0m_n157), .Y(c0sm_b0m_v0m_n45));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u122 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n44), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n150), .C0(c0sm_b0m_v0m_n152), .Y(c0sm_b0m_v0m_n151));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u121 (.A(c0sm_b0m_v0m_n151), .Y(c0sm_b0m_v0m_n42));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u115 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n41), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n144), .C0(c0sm_b0m_v0m_n146), .Y(c0sm_b0m_v0m_n145));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u114 (.A(c0sm_b0m_v0m_n145), .Y(c0sm_b0m_v0m_n39));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u108 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n38), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n138), .C0(c0sm_b0m_v0m_n140), .Y(c0sm_b0m_v0m_n139));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u107 (.A(c0sm_b0m_v0m_n139), .Y(c0sm_b0m_v0m_n36));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u101 (.A0(c0sm_b0m_v0m_n111), .A1(c0sm_b0m_v0m_n35), .B0(c0sm_b0m_v0m_n110), .B1(c0sm_b0m_v0m_n131), .C0(c0sm_b0m_v0m_n133), .Y(c0sm_b0m_v0m_n132));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u100 (.A(c0sm_b0m_v0m_n132), .Y(c0sm_b0m_v0m_n33));
endmodule
module mux21i_oai221_mx38 
(
  c0sm_b0m_v0m_n105, 
  c0sm_b0m_v0m_n110, 
  c0sm_b0m_v0m_n111, 
  c0sm_b0m_v0m_n112, 
  c0sm_b0m_v0m_n122, 
  c0sm_b0m_v0m_n124, 
  c0sm_b0m_v0m_n23, 
  c0sm_b0m_v0m_n29, 
  c0sm_b0m_v0m_n27,
  c0sm_b0m_v0m_n32
);
  input c0sm_b0m_v0m_n105;
  input c0sm_b0m_v0m_n110;
  input c0sm_b0m_v0m_n111;
  input c0sm_b0m_v0m_n112;
  input c0sm_b0m_v0m_n122;
  input c0sm_b0m_v0m_n124;
  input c0sm_b0m_v0m_n23;
  input c0sm_b0m_v0m_n29;
  output c0sm_b0m_v0m_n27;
  output c0sm_b0m_v0m_n32;

  // moduleNum: x38
  // type: mux21i_oai221
  // conflicting modules: 
  // number of bit inputs: 8
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1058/1070
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:245 c0sm_b0m_v0m_n32 c0sm_b0m_v0m_n27 
  // group: sel; nodes: [ c0sm_b0m_v0m_n111 c0sm_b0m_v0m_n110 ]

  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u93 (.A0(c0sm_b0m_v0m_n110), .A1(c0sm_b0m_v0m_n122), .B0(c0sm_b0m_v0m_n111), .B1(c0sm_b0m_v0m_n29), .C0(c0sm_b0m_v0m_n124), .Y(c0sm_b0m_v0m_n32));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u86 (.A0(c0sm_b0m_v0m_n110), .A1(c0sm_b0m_v0m_n105), .B0(c0sm_b0m_v0m_n111), .B1(c0sm_b0m_v0m_n23), .C0(c0sm_b0m_v0m_n112), .Y(c0sm_b0m_v0m_n27));
endmodule
module reg_mx39 
(
  c0nm_b0m_v0m_n11, 
  c0nm_b0m_v0m_n262, 
  c0nm_b0m_v0m_n263, 
  clk, 
  c0nm_b0m_rdata_0_,
  c0nm_b0m_rdata_1_
);
  input c0nm_b0m_v0m_n11;
  input c0nm_b0m_v0m_n262;
  input c0nm_b0m_v0m_n263;
  input clk;
  output c0nm_b0m_rdata_0_;
  output c0nm_b0m_rdata_1_;
  wire c0nm_b0m_v0m_n206;
  wire c0nm_b0m_v0m_n207;

  // moduleNum: x39
  // type: reg
  // conflicting modules: 
  // number of bit inputs: 4
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 6
  // number of non-inferred gates: 0
  // ILP vars: 1071/1073
  // type: INFERRED
  // marked bad? no
  // group: aux; nodes: [ clk ]
  // group: sel; nodes: [ c0nm_b0m_v0m_n11 ]

  MXT2_X0P5M_A12TR c0nm_b0m_v0m_u196 (.A(c0nm_b0m_v0m_n263), .B(c0nm_b0m_rdata_1_), .S0(c0nm_b0m_v0m_n11), .Y(c0nm_b0m_v0m_n206));
  MXT2_X0P5M_A12TR c0nm_b0m_v0m_u194 (.A(c0nm_b0m_v0m_n262), .B(c0nm_b0m_rdata_0_), .S0(c0nm_b0m_v0m_n11), .Y(c0nm_b0m_v0m_n207));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_0_ (.CK(clk), .Q(c0nm_b0m_rdata_0_), .D(c0nm_b0m_v0m_n207));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_1_ (.CK(clk), .Q(c0nm_b0m_rdata_1_), .D(c0nm_b0m_v0m_n206));
endmodule
module reg_mx40 
(
  c0sm_b0m_v0m_n11, 
  c0sm_b0m_v0m_n262, 
  c0sm_b0m_v0m_n263, 
  clk, 
  c0sm_b0m_rdata_0_,
  c0sm_b0m_rdata_1_
);
  input c0sm_b0m_v0m_n11;
  input c0sm_b0m_v0m_n262;
  input c0sm_b0m_v0m_n263;
  input clk;
  output c0sm_b0m_rdata_0_;
  output c0sm_b0m_rdata_1_;
  wire c0sm_b0m_v0m_n331;
  wire c0sm_b0m_v0m_n332;

  // moduleNum: x40
  // type: reg
  // conflicting modules: 
  // number of bit inputs: 4
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 6
  // number of non-inferred gates: 0
  // ILP vars: 1074/1076
  // type: INFERRED
  // marked bad? no
  // group: aux; nodes: [ clk ]
  // group: sel; nodes: [ c0sm_b0m_v0m_n11 ]

  MXT2_X0P5M_A12TR c0sm_b0m_v0m_u196 (.A(c0sm_b0m_v0m_n263), .B(c0sm_b0m_rdata_1_), .S0(c0sm_b0m_v0m_n11), .Y(c0sm_b0m_v0m_n332));
  MXT2_X0P5M_A12TR c0sm_b0m_v0m_u194 (.A(c0sm_b0m_v0m_n262), .B(c0sm_b0m_rdata_0_), .S0(c0sm_b0m_v0m_n11), .Y(c0sm_b0m_v0m_n331));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_0_ (.CK(clk), .Q(c0sm_b0m_rdata_0_), .D(c0sm_b0m_v0m_n331));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_1_ (.CK(clk), .Q(c0sm_b0m_rdata_1_), .D(c0sm_b0m_v0m_n332));
endmodule
module reg_mx41 
(
  c0nm_b0m_v0m_n101, 
  c0nm_b0m_v0m_n97, 
  c0nm_b0m_v0m_n98, 
  clk, 
  c0nm_b0m_v0m_n60,
  c0nm_b0m_v0m_n61
);
  input c0nm_b0m_v0m_n101;
  input c0nm_b0m_v0m_n97;
  input c0nm_b0m_v0m_n98;
  input clk;
  output c0nm_b0m_v0m_n60;
  output c0nm_b0m_v0m_n61;
  wire c0nm_b0m_v0m_n230;
  wire c0nm_b0m_v0m_n231;

  // moduleNum: x41
  // type: reg
  // conflicting modules: 
  // number of bit inputs: 4
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 6
  // number of non-inferred gates: 0
  // ILP vars: 1077/1079
  // type: INFERRED
  // marked bad? no
  // group: aux; nodes: [ clk ]
  // group: sel; nodes: [ c0nm_b0m_v0m_n98 ]

  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u67 (.A(c0nm_b0m_v0m_n60), .B(c0nm_b0m_v0m_n101), .S0(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n230));
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u65 (.A(c0nm_b0m_v0m_n61), .B(c0nm_b0m_v0m_n97), .S0(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n231));
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_0_ (.CK(clk), .QN(c0nm_b0m_v0m_n61), .D(c0nm_b0m_v0m_n231));
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_1_ (.CK(clk), .QN(c0nm_b0m_v0m_n60), .D(c0nm_b0m_v0m_n230));
endmodule
module reg_mx42 
(
  c0sm_b0m_v0m_n101, 
  c0sm_b0m_v0m_n97, 
  c0sm_b0m_v0m_n98, 
  clk, 
  c0sm_b0m_v0m_n343,
  c0sm_b0m_v0m_n344
);
  input c0sm_b0m_v0m_n101;
  input c0sm_b0m_v0m_n97;
  input c0sm_b0m_v0m_n98;
  input clk;
  output c0sm_b0m_v0m_n343;
  output c0sm_b0m_v0m_n344;
  wire c0sm_b0m_v0m_n307;
  wire c0sm_b0m_v0m_n308;

  // moduleNum: x42
  // type: reg
  // conflicting modules: 
  // number of bit inputs: 4
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 6
  // number of non-inferred gates: 0
  // ILP vars: 1080/1082
  // type: INFERRED
  // marked bad? no
  // group: aux; nodes: [ clk ]
  // group: sel; nodes: [ c0sm_b0m_v0m_n98 ]

  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u67 (.A(c0sm_b0m_v0m_n344), .B(c0sm_b0m_v0m_n101), .S0(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n308));
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u65 (.A(c0sm_b0m_v0m_n343), .B(c0sm_b0m_v0m_n97), .S0(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n307));
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_0_ (.CK(clk), .QN(c0sm_b0m_v0m_n343), .D(c0sm_b0m_v0m_n307));
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_1_ (.CK(clk), .QN(c0sm_b0m_v0m_n344), .D(c0sm_b0m_v0m_n308));
endmodule
module reg_mx43 
(
  c0nm_b0m_headflit_10_, 
  c0nm_b0m_headflit_11_, 
  c0nm_b0m_headflit_8_, 
  c0nm_b0m_headflit_9_, 
  c0nm_b0m_v0m_n10, 
  c0nm_b0m_v0m_n11, 
  c0nm_headflit_2_, 
  c0nm_headflit_3_, 
  c0nm_headflit_4_, 
  c0nm_headflit_5_, 
  c0nm_headflit_6_, 
  c0nm_headflit_7_, 
  clk, 
  c0nm_b0m_rdata_10_,
  c0nm_b0m_rdata_11_,
  c0nm_b0m_rdata_2_,
  c0nm_b0m_rdata_3_,
  c0nm_b0m_rdata_4_,
  c0nm_b0m_rdata_5_,
  c0nm_b0m_rdata_6_,
  c0nm_b0m_rdata_7_,
  c0nm_b0m_rdata_8_,
  c0nm_b0m_rdata_9_
);
  input c0nm_b0m_headflit_10_;
  input c0nm_b0m_headflit_11_;
  input c0nm_b0m_headflit_8_;
  input c0nm_b0m_headflit_9_;
  input c0nm_b0m_v0m_n10;
  input c0nm_b0m_v0m_n11;
  input c0nm_headflit_2_;
  input c0nm_headflit_3_;
  input c0nm_headflit_4_;
  input c0nm_headflit_5_;
  input c0nm_headflit_6_;
  input c0nm_headflit_7_;
  input clk;
  output c0nm_b0m_rdata_10_;
  output c0nm_b0m_rdata_11_;
  output c0nm_b0m_rdata_2_;
  output c0nm_b0m_rdata_3_;
  output c0nm_b0m_rdata_4_;
  output c0nm_b0m_rdata_5_;
  output c0nm_b0m_rdata_6_;
  output c0nm_b0m_rdata_7_;
  output c0nm_b0m_rdata_8_;
  output c0nm_b0m_rdata_9_;
  wire c0nm_b0m_v0m_n196;
  wire c0nm_b0m_v0m_n197;
  wire c0nm_b0m_v0m_n198;
  wire c0nm_b0m_v0m_n199;
  wire c0nm_b0m_v0m_n200;
  wire c0nm_b0m_v0m_n201;
  wire c0nm_b0m_v0m_n202;
  wire c0nm_b0m_v0m_n203;
  wire c0nm_b0m_v0m_n204;
  wire c0nm_b0m_v0m_n205;

  // moduleNum: x43
  // type: reg
  // conflicting modules: 
  // number of bit inputs: 13
  // number of bit outputs: 10
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 30
  // number of non-inferred gates: 0
  // ILP vars: 1083/1093
  // type: INFERRED
  // marked bad? no
  // group: aux; nodes: [ clk ]
  // group: sel; nodes: [ c0nm_b0m_v0m_n11 c0nm_b0m_v0m_n10 ]

  AO22_X0P5M_A12TR c0nm_b0m_v0m_u207 (.A0(c0nm_b0m_rdata_11_), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_b0m_headflit_11_), .Y(c0nm_b0m_v0m_n196));
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u206 (.A0(c0nm_b0m_rdata_10_), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_b0m_headflit_10_), .Y(c0nm_b0m_v0m_n197));
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u205 (.A0(c0nm_b0m_rdata_9_), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_b0m_headflit_9_), .Y(c0nm_b0m_v0m_n198));
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u204 (.A0(c0nm_b0m_rdata_8_), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_b0m_headflit_8_), .Y(c0nm_b0m_v0m_n199));
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u203 (.A0(c0nm_b0m_rdata_7_), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit_7_), .Y(c0nm_b0m_v0m_n200));
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u202 (.A0(c0nm_b0m_rdata_6_), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit_6_), .Y(c0nm_b0m_v0m_n201));
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u201 (.A0(c0nm_b0m_rdata_5_), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit_5_), .Y(c0nm_b0m_v0m_n202));
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u200 (.A0(c0nm_b0m_rdata_4_), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit_4_), .Y(c0nm_b0m_v0m_n203));
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u199 (.A0(c0nm_b0m_rdata_3_), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit_3_), .Y(c0nm_b0m_v0m_n204));
  AO22_X0P5M_A12TR c0nm_b0m_v0m_u198 (.A0(c0nm_b0m_rdata_2_), .A1(c0nm_b0m_v0m_n11), .B0(c0nm_b0m_v0m_n10), .B1(c0nm_headflit_2_), .Y(c0nm_b0m_v0m_n205));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_10_ (.CK(clk), .Q(c0nm_b0m_rdata_10_), .D(c0nm_b0m_v0m_n197));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_11_ (.CK(clk), .Q(c0nm_b0m_rdata_11_), .D(c0nm_b0m_v0m_n196));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_2_ (.CK(clk), .Q(c0nm_b0m_rdata_2_), .D(c0nm_b0m_v0m_n205));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_3_ (.CK(clk), .Q(c0nm_b0m_rdata_3_), .D(c0nm_b0m_v0m_n204));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_4_ (.CK(clk), .Q(c0nm_b0m_rdata_4_), .D(c0nm_b0m_v0m_n203));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_5_ (.CK(clk), .Q(c0nm_b0m_rdata_5_), .D(c0nm_b0m_v0m_n202));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_6_ (.CK(clk), .Q(c0nm_b0m_rdata_6_), .D(c0nm_b0m_v0m_n201));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_7_ (.CK(clk), .Q(c0nm_b0m_rdata_7_), .D(c0nm_b0m_v0m_n200));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_8_ (.CK(clk), .Q(c0nm_b0m_rdata_8_), .D(c0nm_b0m_v0m_n199));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_rdata_reg_9_ (.CK(clk), .Q(c0nm_b0m_rdata_9_), .D(c0nm_b0m_v0m_n198));
endmodule
module reg_mx44 
(
  c0sm_b0m_headflit_10_, 
  c0sm_b0m_headflit_11_, 
  c0sm_b0m_headflit_8_, 
  c0sm_b0m_headflit_9_, 
  c0sm_b0m_v0m_n10, 
  c0sm_b0m_v0m_n11, 
  c0sm_headflit_2_, 
  c0sm_headflit_3_, 
  c0sm_headflit_4_, 
  c0sm_headflit_5_, 
  c0sm_headflit_6_, 
  c0sm_headflit_7_, 
  clk, 
  c0sm_b0m_rdata_10_,
  c0sm_b0m_rdata_11_,
  c0sm_b0m_rdata_2_,
  c0sm_b0m_rdata_3_,
  c0sm_b0m_rdata_4_,
  c0sm_b0m_rdata_5_,
  c0sm_b0m_rdata_6_,
  c0sm_b0m_rdata_7_,
  c0sm_b0m_rdata_8_,
  c0sm_b0m_rdata_9_
);
  input c0sm_b0m_headflit_10_;
  input c0sm_b0m_headflit_11_;
  input c0sm_b0m_headflit_8_;
  input c0sm_b0m_headflit_9_;
  input c0sm_b0m_v0m_n10;
  input c0sm_b0m_v0m_n11;
  input c0sm_headflit_2_;
  input c0sm_headflit_3_;
  input c0sm_headflit_4_;
  input c0sm_headflit_5_;
  input c0sm_headflit_6_;
  input c0sm_headflit_7_;
  input clk;
  output c0sm_b0m_rdata_10_;
  output c0sm_b0m_rdata_11_;
  output c0sm_b0m_rdata_2_;
  output c0sm_b0m_rdata_3_;
  output c0sm_b0m_rdata_4_;
  output c0sm_b0m_rdata_5_;
  output c0sm_b0m_rdata_6_;
  output c0sm_b0m_rdata_7_;
  output c0sm_b0m_rdata_8_;
  output c0sm_b0m_rdata_9_;
  wire c0sm_b0m_v0m_n333;
  wire c0sm_b0m_v0m_n334;
  wire c0sm_b0m_v0m_n335;
  wire c0sm_b0m_v0m_n336;
  wire c0sm_b0m_v0m_n337;
  wire c0sm_b0m_v0m_n338;
  wire c0sm_b0m_v0m_n339;
  wire c0sm_b0m_v0m_n340;
  wire c0sm_b0m_v0m_n341;
  wire c0sm_b0m_v0m_n342;

  // moduleNum: x44
  // type: reg
  // conflicting modules: 
  // number of bit inputs: 13
  // number of bit outputs: 10
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 30
  // number of non-inferred gates: 0
  // ILP vars: 1094/1104
  // type: INFERRED
  // marked bad? no
  // group: aux; nodes: [ clk ]
  // group: sel; nodes: [ c0sm_b0m_v0m_n11 c0sm_b0m_v0m_n10 ]

  AO22_X0P5M_A12TR c0sm_b0m_v0m_u207 (.A0(c0sm_b0m_rdata_11_), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_b0m_headflit_11_), .Y(c0sm_b0m_v0m_n342));
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u206 (.A0(c0sm_b0m_rdata_10_), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_b0m_headflit_10_), .Y(c0sm_b0m_v0m_n341));
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u205 (.A0(c0sm_b0m_rdata_9_), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_b0m_headflit_9_), .Y(c0sm_b0m_v0m_n340));
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u204 (.A0(c0sm_b0m_rdata_8_), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_b0m_headflit_8_), .Y(c0sm_b0m_v0m_n339));
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u203 (.A0(c0sm_b0m_rdata_7_), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit_7_), .Y(c0sm_b0m_v0m_n338));
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u202 (.A0(c0sm_b0m_rdata_6_), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit_6_), .Y(c0sm_b0m_v0m_n337));
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u201 (.A0(c0sm_b0m_rdata_5_), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit_5_), .Y(c0sm_b0m_v0m_n336));
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u200 (.A0(c0sm_b0m_rdata_4_), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit_4_), .Y(c0sm_b0m_v0m_n335));
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u199 (.A0(c0sm_b0m_rdata_3_), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit_3_), .Y(c0sm_b0m_v0m_n334));
  AO22_X0P5M_A12TR c0sm_b0m_v0m_u198 (.A0(c0sm_b0m_rdata_2_), .A1(c0sm_b0m_v0m_n11), .B0(c0sm_b0m_v0m_n10), .B1(c0sm_headflit_2_), .Y(c0sm_b0m_v0m_n333));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_10_ (.CK(clk), .Q(c0sm_b0m_rdata_10_), .D(c0sm_b0m_v0m_n341));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_11_ (.CK(clk), .Q(c0sm_b0m_rdata_11_), .D(c0sm_b0m_v0m_n342));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_2_ (.CK(clk), .Q(c0sm_b0m_rdata_2_), .D(c0sm_b0m_v0m_n333));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_3_ (.CK(clk), .Q(c0sm_b0m_rdata_3_), .D(c0sm_b0m_v0m_n334));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_4_ (.CK(clk), .Q(c0sm_b0m_rdata_4_), .D(c0sm_b0m_v0m_n335));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_5_ (.CK(clk), .Q(c0sm_b0m_rdata_5_), .D(c0sm_b0m_v0m_n336));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_6_ (.CK(clk), .Q(c0sm_b0m_rdata_6_), .D(c0sm_b0m_v0m_n337));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_7_ (.CK(clk), .Q(c0sm_b0m_rdata_7_), .D(c0sm_b0m_v0m_n338));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_8_ (.CK(clk), .Q(c0sm_b0m_rdata_8_), .D(c0sm_b0m_v0m_n339));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_rdata_reg_9_ (.CK(clk), .Q(c0sm_b0m_rdata_9_), .D(c0sm_b0m_v0m_n340));
endmodule
module reg_mx45 
(
  c0nm_b0m_v0m_n102, 
  c0nm_b0m_v0m_n103, 
  c0nm_b0m_v0m_n17, 
  c0nm_b0m_v0m_n19, 
  c0nm_b0m_v0m_n33, 
  c0nm_b0m_v0m_n34, 
  c0nm_b0m_v0m_n36, 
  c0nm_b0m_v0m_n37, 
  c0nm_b0m_v0m_n39, 
  c0nm_b0m_v0m_n40, 
  c0nm_b0m_v0m_n42, 
  c0nm_b0m_v0m_n43, 
  c0nm_b0m_v0m_n45, 
  c0nm_b0m_v0m_n46, 
  c0nm_b0m_v0m_n48, 
  c0nm_b0m_v0m_n49, 
  c0nm_b0m_v0m_n63, 
  c0nm_b0m_v0m_n64, 
  c0nm_b0m_v0m_n66, 
  c0nm_b0m_v0m_n67, 
  c0nm_b0m_v0m_n69, 
  c0nm_b0m_v0m_n70, 
  c0nm_b0m_v0m_n98, 
  clk, 
  c0nm_b0m_v0m_n50,
  c0nm_b0m_v0m_n51,
  c0nm_b0m_v0m_n52,
  c0nm_b0m_v0m_n53,
  c0nm_b0m_v0m_n54,
  c0nm_b0m_v0m_n55,
  c0nm_b0m_v0m_n56,
  c0nm_b0m_v0m_n57,
  c0nm_b0m_v0m_n58,
  c0nm_b0m_v0m_n59
);
  input c0nm_b0m_v0m_n102;
  input c0nm_b0m_v0m_n103;
  input c0nm_b0m_v0m_n17;
  input c0nm_b0m_v0m_n19;
  input c0nm_b0m_v0m_n33;
  input c0nm_b0m_v0m_n34;
  input c0nm_b0m_v0m_n36;
  input c0nm_b0m_v0m_n37;
  input c0nm_b0m_v0m_n39;
  input c0nm_b0m_v0m_n40;
  input c0nm_b0m_v0m_n42;
  input c0nm_b0m_v0m_n43;
  input c0nm_b0m_v0m_n45;
  input c0nm_b0m_v0m_n46;
  input c0nm_b0m_v0m_n48;
  input c0nm_b0m_v0m_n49;
  input c0nm_b0m_v0m_n63;
  input c0nm_b0m_v0m_n64;
  input c0nm_b0m_v0m_n66;
  input c0nm_b0m_v0m_n67;
  input c0nm_b0m_v0m_n69;
  input c0nm_b0m_v0m_n70;
  input c0nm_b0m_v0m_n98;
  input clk;
  output c0nm_b0m_v0m_n50;
  output c0nm_b0m_v0m_n51;
  output c0nm_b0m_v0m_n52;
  output c0nm_b0m_v0m_n53;
  output c0nm_b0m_v0m_n54;
  output c0nm_b0m_v0m_n55;
  output c0nm_b0m_v0m_n56;
  output c0nm_b0m_v0m_n57;
  output c0nm_b0m_v0m_n58;
  output c0nm_b0m_v0m_n59;
  wire c0nm_b0m_v0m_n220;
  wire c0nm_b0m_v0m_n221;
  wire c0nm_b0m_v0m_n222;
  wire c0nm_b0m_v0m_n223;
  wire c0nm_b0m_v0m_n224;
  wire c0nm_b0m_v0m_n225;
  wire c0nm_b0m_v0m_n226;
  wire c0nm_b0m_v0m_n227;
  wire c0nm_b0m_v0m_n228;
  wire c0nm_b0m_v0m_n229;

  // moduleNum: x45
  // type: reg
  // conflicting modules: 
  // number of bit inputs: 24
  // number of bit outputs: 10
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 30
  // number of non-inferred gates: 0
  // ILP vars: 1105/1115
  // type: INFERRED
  // marked bad? no
  // group: aux; nodes: [ clk ]
  // group: sel; nodes: [ c0nm_b0m_v0m_n102 c0nm_b0m_v0m_n98 c0nm_b0m_v0m_n103 ]

  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u78 (.A0(c0nm_b0m_v0m_n19), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n17), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n50), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n220));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u77 (.A0(c0nm_b0m_v0m_n70), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n69), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n51), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n221));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u76 (.A0(c0nm_b0m_v0m_n67), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n66), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n52), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n222));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u75 (.A0(c0nm_b0m_v0m_n64), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n63), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n53), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n223));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u74 (.A0(c0nm_b0m_v0m_n49), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n48), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n54), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n224));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u73 (.A0(c0nm_b0m_v0m_n46), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n45), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n55), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n225));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u72 (.A0(c0nm_b0m_v0m_n43), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n42), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n56), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n226));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u71 (.A0(c0nm_b0m_v0m_n40), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n39), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n57), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n227));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u70 (.A0(c0nm_b0m_v0m_n37), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n36), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n58), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n228));
  OAI222_X0P5M_A12TR c0nm_b0m_v0m_u69 (.A0(c0nm_b0m_v0m_n34), .A1(c0nm_b0m_v0m_n102), .B0(c0nm_b0m_v0m_n33), .B1(c0nm_b0m_v0m_n103), .C0(c0nm_b0m_v0m_n59), .C1(c0nm_b0m_v0m_n98), .Y(c0nm_b0m_v0m_n229));
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_2_ (.CK(clk), .QN(c0nm_b0m_v0m_n59), .D(c0nm_b0m_v0m_n229));
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_3_ (.CK(clk), .QN(c0nm_b0m_v0m_n58), .D(c0nm_b0m_v0m_n228));
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_4_ (.CK(clk), .QN(c0nm_b0m_v0m_n57), .D(c0nm_b0m_v0m_n227));
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_5_ (.CK(clk), .QN(c0nm_b0m_v0m_n56), .D(c0nm_b0m_v0m_n226));
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_6_ (.CK(clk), .QN(c0nm_b0m_v0m_n55), .D(c0nm_b0m_v0m_n225));
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_7_ (.CK(clk), .QN(c0nm_b0m_v0m_n54), .D(c0nm_b0m_v0m_n224));
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_8_ (.CK(clk), .QN(c0nm_b0m_v0m_n53), .D(c0nm_b0m_v0m_n223));
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_9_ (.CK(clk), .QN(c0nm_b0m_v0m_n52), .D(c0nm_b0m_v0m_n222));
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_10_ (.CK(clk), .QN(c0nm_b0m_v0m_n51), .D(c0nm_b0m_v0m_n221));
  DFFQN_X1M_A12TR c0nm_b0m_v0m_buffers1_reg_11_ (.CK(clk), .QN(c0nm_b0m_v0m_n50), .D(c0nm_b0m_v0m_n220));
endmodule
module reg_mx46 
(
  c0sm_b0m_v0m_n102, 
  c0sm_b0m_v0m_n103, 
  c0sm_b0m_v0m_n17, 
  c0sm_b0m_v0m_n19, 
  c0sm_b0m_v0m_n33, 
  c0sm_b0m_v0m_n34, 
  c0sm_b0m_v0m_n36, 
  c0sm_b0m_v0m_n37, 
  c0sm_b0m_v0m_n39, 
  c0sm_b0m_v0m_n40, 
  c0sm_b0m_v0m_n42, 
  c0sm_b0m_v0m_n43, 
  c0sm_b0m_v0m_n45, 
  c0sm_b0m_v0m_n46, 
  c0sm_b0m_v0m_n48, 
  c0sm_b0m_v0m_n49, 
  c0sm_b0m_v0m_n63, 
  c0sm_b0m_v0m_n64, 
  c0sm_b0m_v0m_n66, 
  c0sm_b0m_v0m_n67, 
  c0sm_b0m_v0m_n69, 
  c0sm_b0m_v0m_n70, 
  c0sm_b0m_v0m_n98, 
  clk, 
  c0sm_b0m_v0m_n345,
  c0sm_b0m_v0m_n346,
  c0sm_b0m_v0m_n347,
  c0sm_b0m_v0m_n348,
  c0sm_b0m_v0m_n349,
  c0sm_b0m_v0m_n350,
  c0sm_b0m_v0m_n351,
  c0sm_b0m_v0m_n352,
  c0sm_b0m_v0m_n353,
  c0sm_b0m_v0m_n354
);
  input c0sm_b0m_v0m_n102;
  input c0sm_b0m_v0m_n103;
  input c0sm_b0m_v0m_n17;
  input c0sm_b0m_v0m_n19;
  input c0sm_b0m_v0m_n33;
  input c0sm_b0m_v0m_n34;
  input c0sm_b0m_v0m_n36;
  input c0sm_b0m_v0m_n37;
  input c0sm_b0m_v0m_n39;
  input c0sm_b0m_v0m_n40;
  input c0sm_b0m_v0m_n42;
  input c0sm_b0m_v0m_n43;
  input c0sm_b0m_v0m_n45;
  input c0sm_b0m_v0m_n46;
  input c0sm_b0m_v0m_n48;
  input c0sm_b0m_v0m_n49;
  input c0sm_b0m_v0m_n63;
  input c0sm_b0m_v0m_n64;
  input c0sm_b0m_v0m_n66;
  input c0sm_b0m_v0m_n67;
  input c0sm_b0m_v0m_n69;
  input c0sm_b0m_v0m_n70;
  input c0sm_b0m_v0m_n98;
  input clk;
  output c0sm_b0m_v0m_n345;
  output c0sm_b0m_v0m_n346;
  output c0sm_b0m_v0m_n347;
  output c0sm_b0m_v0m_n348;
  output c0sm_b0m_v0m_n349;
  output c0sm_b0m_v0m_n350;
  output c0sm_b0m_v0m_n351;
  output c0sm_b0m_v0m_n352;
  output c0sm_b0m_v0m_n353;
  output c0sm_b0m_v0m_n354;
  wire c0sm_b0m_v0m_n309;
  wire c0sm_b0m_v0m_n310;
  wire c0sm_b0m_v0m_n311;
  wire c0sm_b0m_v0m_n312;
  wire c0sm_b0m_v0m_n313;
  wire c0sm_b0m_v0m_n314;
  wire c0sm_b0m_v0m_n315;
  wire c0sm_b0m_v0m_n316;
  wire c0sm_b0m_v0m_n317;
  wire c0sm_b0m_v0m_n318;

  // moduleNum: x46
  // type: reg
  // conflicting modules: 
  // number of bit inputs: 24
  // number of bit outputs: 10
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 30
  // number of non-inferred gates: 0
  // ILP vars: 1116/1126
  // type: INFERRED
  // marked bad? no
  // group: aux; nodes: [ clk ]
  // group: sel; nodes: [ c0sm_b0m_v0m_n102 c0sm_b0m_v0m_n98 c0sm_b0m_v0m_n103 ]

  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u78 (.A0(c0sm_b0m_v0m_n19), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n17), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n354), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n318));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u77 (.A0(c0sm_b0m_v0m_n70), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n69), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n353), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n317));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u76 (.A0(c0sm_b0m_v0m_n67), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n66), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n352), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n316));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u75 (.A0(c0sm_b0m_v0m_n64), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n63), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n351), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n315));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u74 (.A0(c0sm_b0m_v0m_n49), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n48), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n350), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n314));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u73 (.A0(c0sm_b0m_v0m_n46), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n45), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n349), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n313));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u72 (.A0(c0sm_b0m_v0m_n43), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n42), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n348), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n312));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u71 (.A0(c0sm_b0m_v0m_n40), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n39), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n347), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n311));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u70 (.A0(c0sm_b0m_v0m_n37), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n36), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n346), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n310));
  OAI222_X0P5M_A12TR c0sm_b0m_v0m_u69 (.A0(c0sm_b0m_v0m_n34), .A1(c0sm_b0m_v0m_n102), .B0(c0sm_b0m_v0m_n33), .B1(c0sm_b0m_v0m_n103), .C0(c0sm_b0m_v0m_n345), .C1(c0sm_b0m_v0m_n98), .Y(c0sm_b0m_v0m_n309));
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_2_ (.CK(clk), .QN(c0sm_b0m_v0m_n345), .D(c0sm_b0m_v0m_n309));
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_3_ (.CK(clk), .QN(c0sm_b0m_v0m_n346), .D(c0sm_b0m_v0m_n310));
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_4_ (.CK(clk), .QN(c0sm_b0m_v0m_n347), .D(c0sm_b0m_v0m_n311));
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_5_ (.CK(clk), .QN(c0sm_b0m_v0m_n348), .D(c0sm_b0m_v0m_n312));
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_6_ (.CK(clk), .QN(c0sm_b0m_v0m_n349), .D(c0sm_b0m_v0m_n313));
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_7_ (.CK(clk), .QN(c0sm_b0m_v0m_n350), .D(c0sm_b0m_v0m_n314));
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_8_ (.CK(clk), .QN(c0sm_b0m_v0m_n351), .D(c0sm_b0m_v0m_n315));
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_9_ (.CK(clk), .QN(c0sm_b0m_v0m_n352), .D(c0sm_b0m_v0m_n316));
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_10_ (.CK(clk), .QN(c0sm_b0m_v0m_n353), .D(c0sm_b0m_v0m_n317));
  DFFQN_X1M_A12TR c0sm_b0m_v0m_buffers1_reg_11_ (.CK(clk), .QN(c0sm_b0m_v0m_n354), .D(c0sm_b0m_v0m_n318));
endmodule
module decoder24_mx47 
(
  swalloc_resp_0_0_, 
  swalloc_resp_1_0_, 
  colsel0_0_,
  colsel0_1_
);
  input swalloc_resp_0_0_;
  input swalloc_resp_1_0_;
  output colsel0_0_;
  output colsel0_1_;

  // moduleNum: x47
  // type: decoder24
  // conflicting modules: 
  // number of bit inputs: 2
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1135/1135
  // type: INFERRED
  // marked bad? no
  // group: sel; nodes: [ swalloc_resp_0[0] swalloc_resp_1[0] ]

  NAND2B_X0P5M_A12TR d0m_u2 (.AN(swalloc_resp_1_0_), .B(swalloc_resp_0_0_), .Y(colsel0_0_));
  NOR2_X0P5A_A12TR d0m_u1 (.A(swalloc_resp_1_0_), .B(swalloc_resp_0_0_), .Y(colsel0_1_));
endmodule
module decoder24_mx48 
(
  swalloc_resp_0_1_, 
  swalloc_resp_1_1_, 
  colsel1_0_,
  colsel1_1_
);
  input swalloc_resp_0_1_;
  input swalloc_resp_1_1_;
  output colsel1_0_;
  output colsel1_1_;

  // moduleNum: x48
  // type: decoder24
  // conflicting modules: 
  // number of bit inputs: 2
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1136/1136
  // type: INFERRED
  // marked bad? no
  // group: sel; nodes: [ swalloc_resp_0[1] swalloc_resp_1[1] ]

  NAND2B_X0P5M_A12TR d1m_u2 (.AN(swalloc_resp_1_1_), .B(swalloc_resp_0_1_), .Y(colsel1_0_));
  NOR2_X0P5A_A12TR d1m_u1 (.A(swalloc_resp_1_1_), .B(swalloc_resp_0_1_), .Y(colsel1_1_));
endmodule
module decoder24_mx49 
(
  s0m_o0nm_state_credits_0_, 
  s0m_o0nm_state_credits_1_, 
  s0m_o0nm_n18,
  s0m_o0nm_n22
);
  input s0m_o0nm_state_credits_0_;
  input s0m_o0nm_state_credits_1_;
  output s0m_o0nm_n18;
  output s0m_o0nm_n22;

  // moduleNum: x49
  // type: decoder24
  // conflicting modules: 
  // number of bit inputs: 2
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1137/1137
  // type: INFERRED
  // marked bad? no
  // group: sel; nodes: [ s0m_o0nm_state_credits_0_ s0m_o0nm_state_credits_1_ ]

  OR2_X0P5M_A12TR s0m_o0nm_u29 (.A(s0m_o0nm_state_credits_1_), .B(s0m_o0nm_state_credits_0_), .Y(s0m_o0nm_n22));
  NAND2_X0P5A_A12TR s0m_o0nm_u22 (.A(s0m_o0nm_state_credits_1_), .B(s0m_o0nm_state_credits_0_), .Y(s0m_o0nm_n18));
endmodule
module decoder24_mx50 
(
  s0m_o0sm_state_credits_0_, 
  s0m_o0sm_state_credits_1_, 
  s0m_o0sm_n18,
  s0m_o0sm_n22
);
  input s0m_o0sm_state_credits_0_;
  input s0m_o0sm_state_credits_1_;
  output s0m_o0sm_n18;
  output s0m_o0sm_n22;

  // moduleNum: x50
  // type: decoder24
  // conflicting modules: 
  // number of bit inputs: 2
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1138/1138
  // type: INFERRED
  // marked bad? no
  // group: sel; nodes: [ s0m_o0sm_state_credits_0_ s0m_o0sm_state_credits_1_ ]

  OR2_X0P5M_A12TR s0m_o0sm_u29 (.A(s0m_o0sm_state_credits_1_), .B(s0m_o0sm_state_credits_0_), .Y(s0m_o0sm_n22));
  NAND2_X0P5A_A12TR s0m_o0sm_u22 (.A(s0m_o0sm_state_credits_1_), .B(s0m_o0sm_state_credits_0_), .Y(s0m_o0sm_n18));
endmodule
module decoder38_mx51 
(
  creditin_0, 
  s0m_o0nm_n12, 
  s0m_o0nm_n9, 
  s0m_o0nm_n20,
  s0m_o0nm_n6
);
  input creditin_0;
  input s0m_o0nm_n12;
  input s0m_o0nm_n9;
  output s0m_o0nm_n20;
  output s0m_o0nm_n6;
  wire s0m_o0nm_n11;

  // moduleNum: x51
  // type: decoder38
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 3
  // number of non-inferred gates: 0
  // ILP vars: 1147/1147
  // type: INFERRED
  // marked bad? no
  // group: sel; nodes: [ creditin_0 s0m_o0nm_n9 s0m_o0nm_n12 ]

  NOR3_X0P5A_A12TR s0m_o0nm_u27 (.A(s0m_o0nm_n9), .B(creditin_0), .C(s0m_o0nm_n12), .Y(s0m_o0nm_n20));
  INV_X0P5B_A12TR s0m_o0nm_u13 (.A(s0m_o0nm_n12), .Y(s0m_o0nm_n11));
  NOR3_X0P5A_A12TR s0m_o0nm_u12 (.A(s0m_o0nm_n11), .B(creditin_0), .C(s0m_o0nm_n9), .Y(s0m_o0nm_n6));
endmodule
module decoder38_mx52 
(
  creditin_1, 
  s0m_o0sm_n12, 
  s0m_o0sm_n9, 
  s0m_o0sm_n20,
  s0m_o0sm_n6
);
  input creditin_1;
  input s0m_o0sm_n12;
  input s0m_o0sm_n9;
  output s0m_o0sm_n20;
  output s0m_o0sm_n6;
  wire s0m_o0sm_n11;

  // moduleNum: x52
  // type: decoder38
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 3
  // number of non-inferred gates: 0
  // ILP vars: 1148/1148
  // type: INFERRED
  // marked bad? no
  // group: sel; nodes: [ creditin_1 s0m_o0sm_n9 s0m_o0sm_n12 ]

  NOR3_X0P5A_A12TR s0m_o0sm_u27 (.A(s0m_o0sm_n9), .B(creditin_1), .C(s0m_o0sm_n12), .Y(s0m_o0sm_n20));
  INV_X0P5B_A12TR s0m_o0sm_u13 (.A(s0m_o0sm_n12), .Y(s0m_o0sm_n11));
  NOR3_X0P5A_A12TR s0m_o0sm_u12 (.A(s0m_o0sm_n11), .B(creditin_1), .C(s0m_o0sm_n9), .Y(s0m_o0sm_n6));
endmodule
module decoder38_mx53 
(
  c0nm_b0m_v0m_n9, 
  c0nm_b0m_v0m_tail_0_, 
  c0nm_b0m_v0m_tail_1_, 
  c0nm_b0m_v0m_n100,
  c0nm_b0m_v0m_n109,
  c0nm_b0m_v0m_n78,
  c0nm_b0m_v0m_n93,
  c0nm_b0m_v0m_n94,
  c0nm_b0m_v0m_n95
);
  input c0nm_b0m_v0m_n9;
  input c0nm_b0m_v0m_tail_0_;
  input c0nm_b0m_v0m_tail_1_;
  output c0nm_b0m_v0m_n100;
  output c0nm_b0m_v0m_n109;
  output c0nm_b0m_v0m_n78;
  output c0nm_b0m_v0m_n93;
  output c0nm_b0m_v0m_n94;
  output c0nm_b0m_v0m_n95;
  wire c0nm_b0m_v0m_n26;
  wire c0nm_b0m_v0m_n3;
  wire c0nm_b0m_v0m_n7;
  wire c0nm_b0m_v0m_n72;

  // moduleNum: x53
  // type: decoder38
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 6
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 1165/1174
  // type: INFERRED
  // marked bad? no
  // group: sel; nodes: [ c0nm_b0m_v0m_n9 c0nm_b0m_v0m_tail_0_ c0nm_b0m_v0m_tail_1_ ]

  INV_X0P5B_A12TR c0nm_b0m_v0m_u193 (.A(c0nm_b0m_v0m_tail_1_), .Y(c0nm_b0m_v0m_n7));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u192 (.A(c0nm_b0m_v0m_tail_0_), .B(c0nm_b0m_v0m_n7), .C(c0nm_b0m_v0m_n9), .Y(c0nm_b0m_v0m_n93));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u189 (.A(c0nm_b0m_v0m_tail_0_), .Y(c0nm_b0m_v0m_n3));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u188 (.A(c0nm_b0m_v0m_tail_1_), .B(c0nm_b0m_v0m_n3), .C(c0nm_b0m_v0m_n9), .Y(c0nm_b0m_v0m_n94));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u186 (.A(c0nm_b0m_v0m_n3), .B(c0nm_b0m_v0m_n7), .C(c0nm_b0m_v0m_n9), .Y(c0nm_b0m_v0m_n95));
  OAI21_X0P5M_A12TR c0nm_b0m_v0m_u166 (.A0(c0nm_b0m_v0m_n3), .A1(c0nm_b0m_v0m_n7), .B0(c0nm_b0m_v0m_n9), .Y(c0nm_b0m_v0m_n26));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u165 (.A(c0nm_b0m_v0m_n26), .Y(c0nm_b0m_v0m_n72));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u164 (.A(c0nm_b0m_v0m_n93), .B(c0nm_b0m_v0m_n95), .C(c0nm_b0m_v0m_n72), .Y(c0nm_b0m_v0m_n109));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u80 (.A(c0nm_b0m_v0m_n95), .B(c0nm_b0m_v0m_n94), .C(c0nm_b0m_v0m_n72), .Y(c0nm_b0m_v0m_n100));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u61 (.A(c0nm_b0m_v0m_n93), .B(c0nm_b0m_v0m_n94), .C(c0nm_b0m_v0m_n72), .Y(c0nm_b0m_v0m_n78));
endmodule
module decoder38_mx54 
(
  c0sm_b0m_v0m_n355, 
  c0sm_b0m_v0m_tail_0_, 
  c0sm_b0m_v0m_tail_1_, 
  c0sm_b0m_v0m_n100,
  c0sm_b0m_v0m_n109,
  c0sm_b0m_v0m_n78,
  c0sm_b0m_v0m_n93,
  c0sm_b0m_v0m_n94,
  c0sm_b0m_v0m_n95
);
  input c0sm_b0m_v0m_n355;
  input c0sm_b0m_v0m_tail_0_;
  input c0sm_b0m_v0m_tail_1_;
  output c0sm_b0m_v0m_n100;
  output c0sm_b0m_v0m_n109;
  output c0sm_b0m_v0m_n78;
  output c0sm_b0m_v0m_n93;
  output c0sm_b0m_v0m_n94;
  output c0sm_b0m_v0m_n95;
  wire c0sm_b0m_v0m_n26;
  wire c0sm_b0m_v0m_n3;
  wire c0sm_b0m_v0m_n7;
  wire c0sm_b0m_v0m_n72;

  // moduleNum: x54
  // type: decoder38
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 6
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 1197/1206
  // type: INFERRED
  // marked bad? no
  // group: sel; nodes: [ c0sm_b0m_v0m_n355 c0sm_b0m_v0m_tail_0_ c0sm_b0m_v0m_tail_1_ ]

  INV_X0P5B_A12TR c0sm_b0m_v0m_u193 (.A(c0sm_b0m_v0m_tail_1_), .Y(c0sm_b0m_v0m_n7));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u192 (.A(c0sm_b0m_v0m_tail_0_), .B(c0sm_b0m_v0m_n7), .C(c0sm_b0m_v0m_n355), .Y(c0sm_b0m_v0m_n93));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u189 (.A(c0sm_b0m_v0m_tail_0_), .Y(c0sm_b0m_v0m_n3));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u188 (.A(c0sm_b0m_v0m_tail_1_), .B(c0sm_b0m_v0m_n3), .C(c0sm_b0m_v0m_n355), .Y(c0sm_b0m_v0m_n94));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u186 (.A(c0sm_b0m_v0m_n3), .B(c0sm_b0m_v0m_n7), .C(c0sm_b0m_v0m_n355), .Y(c0sm_b0m_v0m_n95));
  OAI21_X0P5M_A12TR c0sm_b0m_v0m_u166 (.A0(c0sm_b0m_v0m_n3), .A1(c0sm_b0m_v0m_n7), .B0(c0sm_b0m_v0m_n355), .Y(c0sm_b0m_v0m_n26));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u165 (.A(c0sm_b0m_v0m_n26), .Y(c0sm_b0m_v0m_n72));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u164 (.A(c0sm_b0m_v0m_n93), .B(c0sm_b0m_v0m_n95), .C(c0sm_b0m_v0m_n72), .Y(c0sm_b0m_v0m_n109));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u80 (.A(c0sm_b0m_v0m_n95), .B(c0sm_b0m_v0m_n94), .C(c0sm_b0m_v0m_n72), .Y(c0sm_b0m_v0m_n100));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u61 (.A(c0sm_b0m_v0m_n93), .B(c0sm_b0m_v0m_n94), .C(c0sm_b0m_v0m_n72), .Y(c0sm_b0m_v0m_n78));
endmodule
module decoder416_mx55 
(
  c0nm_b0m_v0m_head_0_, 
  c0nm_b0m_v0m_head_1_, 
  c0nm_b0m_v0m_head_2_, 
  debitout_0, 
  c0nm_b0m_v0m_n110,
  c0nm_b0m_v0m_n113,
  c0nm_b0m_v0m_n115
);
  input c0nm_b0m_v0m_head_0_;
  input c0nm_b0m_v0m_head_1_;
  input c0nm_b0m_v0m_head_2_;
  input debitout_0;
  output c0nm_b0m_v0m_n110;
  output c0nm_b0m_v0m_n113;
  output c0nm_b0m_v0m_n115;
  wire c0nm_b0m_v0m_n104;
  wire c0nm_b0m_v0m_n15;
  wire c0nm_b0m_v0m_n16;
  wire c0nm_b0m_v0m_n187;
  wire c0nm_b0m_v0m_n192;
  wire c0nm_b0m_v0m_n193;
  wire c0nm_b0m_v0m_n96;

  // moduleNum: x55
  // type: decoder416
  // conflicting modules: 
  // number of bit inputs: 4
  // number of bit outputs: 3
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 1295/1298
  // type: INFERRED
  // marked bad? no
  // group: sel; nodes: [ c0nm_b0m_v0m_head_1_ c0nm_b0m_v0m_head_0_ c0nm_b0m_v0m_head_2_ debitout_0 ]

  INV_X0P5B_A12TR c0nm_b0m_v0m_u278 (.A(c0nm_b0m_v0m_head_0_), .Y(c0nm_b0m_v0m_n16));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u277 (.A(c0nm_b0m_v0m_head_2_), .Y(c0nm_b0m_v0m_n15));
  NAND3_X0P5A_A12TR c0nm_b0m_v0m_u276 (.A(c0nm_b0m_v0m_n16), .B(c0nm_b0m_v0m_n15), .C(c0nm_b0m_v0m_head_1_), .Y(c0nm_b0m_v0m_n187));
  NOR3_X0P5A_A12TR c0nm_b0m_v0m_u272 (.A(c0nm_b0m_v0m_head_1_), .B(c0nm_b0m_v0m_head_2_), .C(c0nm_b0m_v0m_head_0_), .Y(c0nm_b0m_v0m_n193));
  NOR3_X0P5A_A12TR c0nm_b0m_v0m_u271 (.A(c0nm_b0m_v0m_head_1_), .B(c0nm_b0m_v0m_head_2_), .C(c0nm_b0m_v0m_n16), .Y(c0nm_b0m_v0m_n192));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u177 (.A(c0nm_b0m_v0m_n193), .Y(c0nm_b0m_v0m_n96));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u176 (.A(c0nm_b0m_v0m_n192), .Y(c0nm_b0m_v0m_n104));
  OR2_X0P5M_A12TR c0nm_b0m_v0m_u173 (.A(c0nm_b0m_v0m_n187), .B(debitout_0), .Y(c0nm_b0m_v0m_n110));
  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u172 (.A(c0nm_b0m_v0m_n96), .B(debitout_0), .Y(c0nm_b0m_v0m_n115));
  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u171 (.A(c0nm_b0m_v0m_n104), .B(debitout_0), .Y(c0nm_b0m_v0m_n113));
endmodule
module decoder416_mx56 
(
  c0sm_b0m_v0m_head_0_, 
  c0sm_b0m_v0m_head_1_, 
  c0sm_b0m_v0m_head_2_, 
  debitout_1, 
  c0sm_b0m_v0m_n110,
  c0sm_b0m_v0m_n113,
  c0sm_b0m_v0m_n115
);
  input c0sm_b0m_v0m_head_0_;
  input c0sm_b0m_v0m_head_1_;
  input c0sm_b0m_v0m_head_2_;
  input debitout_1;
  output c0sm_b0m_v0m_n110;
  output c0sm_b0m_v0m_n113;
  output c0sm_b0m_v0m_n115;
  wire c0sm_b0m_v0m_n104;
  wire c0sm_b0m_v0m_n15;
  wire c0sm_b0m_v0m_n16;
  wire c0sm_b0m_v0m_n187;
  wire c0sm_b0m_v0m_n192;
  wire c0sm_b0m_v0m_n193;
  wire c0sm_b0m_v0m_n96;

  // moduleNum: x56
  // type: decoder416
  // conflicting modules: 
  // number of bit inputs: 4
  // number of bit outputs: 3
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 1321/1324
  // type: INFERRED
  // marked bad? no
  // group: sel; nodes: [ c0sm_b0m_v0m_head_1_ c0sm_b0m_v0m_head_0_ c0sm_b0m_v0m_head_2_ debitout_1 ]

  INV_X0P5B_A12TR c0sm_b0m_v0m_u278 (.A(c0sm_b0m_v0m_head_0_), .Y(c0sm_b0m_v0m_n16));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u277 (.A(c0sm_b0m_v0m_head_2_), .Y(c0sm_b0m_v0m_n15));
  NAND3_X0P5A_A12TR c0sm_b0m_v0m_u276 (.A(c0sm_b0m_v0m_n16), .B(c0sm_b0m_v0m_n15), .C(c0sm_b0m_v0m_head_1_), .Y(c0sm_b0m_v0m_n187));
  NOR3_X0P5A_A12TR c0sm_b0m_v0m_u272 (.A(c0sm_b0m_v0m_head_1_), .B(c0sm_b0m_v0m_head_2_), .C(c0sm_b0m_v0m_head_0_), .Y(c0sm_b0m_v0m_n193));
  NOR3_X0P5A_A12TR c0sm_b0m_v0m_u271 (.A(c0sm_b0m_v0m_head_1_), .B(c0sm_b0m_v0m_head_2_), .C(c0sm_b0m_v0m_n16), .Y(c0sm_b0m_v0m_n192));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u177 (.A(c0sm_b0m_v0m_n193), .Y(c0sm_b0m_v0m_n96));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u176 (.A(c0sm_b0m_v0m_n192), .Y(c0sm_b0m_v0m_n104));
  OR2_X0P5M_A12TR c0sm_b0m_v0m_u173 (.A(c0sm_b0m_v0m_n187), .B(debitout_1), .Y(c0sm_b0m_v0m_n110));
  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u172 (.A(c0sm_b0m_v0m_n96), .B(debitout_1), .Y(c0sm_b0m_v0m_n115));
  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u171 (.A(c0sm_b0m_v0m_n104), .B(debitout_1), .Y(c0sm_b0m_v0m_n113));
endmodule
module and2gate_mx57 
(
  c0nm_r0m_n15, 
  c0sm_r0m_n15, 
  currx_1_, 
  c0nm_r0m_n16,
  c0sm_r0m_n16
);
  input c0nm_r0m_n15;
  input c0sm_r0m_n15;
  input currx_1_;
  output c0nm_r0m_n16;
  output c0sm_r0m_n16;

  // moduleNum: x57
  // type: and2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1335/1335
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:196 c0sm_r0m_n16 c0nm_r0m_n16 
  // group: sel; nodes: [ currx[1] ]

  AND2_X0P5M_A12TR c0nm_r0m_u16 (.A(c0nm_r0m_n15), .B(currx_1_), .Y(c0nm_r0m_n16));
  AND2_X0P5M_A12TR c0sm_r0m_u16 (.A(c0sm_r0m_n15), .B(currx_1_), .Y(c0sm_r0m_n16));
endmodule
module and2gate_mx58 
(
  c0nm_b0m_n1, 
  flitin_0_10_, 
  flitin_0_11_, 
  flitin_0_2_, 
  flitin_0_3_, 
  flitin_0_4_, 
  flitin_0_5_, 
  flitin_0_6_, 
  flitin_0_7_, 
  flitin_0_8_, 
  flitin_0_9_, 
  c0nm_b0m_wdata_10_,
  c0nm_b0m_wdata_11_,
  c0nm_b0m_wdata_2_,
  c0nm_b0m_wdata_3_,
  c0nm_b0m_wdata_4_,
  c0nm_b0m_wdata_5_,
  c0nm_b0m_wdata_6_,
  c0nm_b0m_wdata_7_,
  c0nm_b0m_wdata_8_,
  c0nm_b0m_wdata_9_
);
  input c0nm_b0m_n1;
  input flitin_0_10_;
  input flitin_0_11_;
  input flitin_0_2_;
  input flitin_0_3_;
  input flitin_0_4_;
  input flitin_0_5_;
  input flitin_0_6_;
  input flitin_0_7_;
  input flitin_0_8_;
  input flitin_0_9_;
  output c0nm_b0m_wdata_10_;
  output c0nm_b0m_wdata_11_;
  output c0nm_b0m_wdata_2_;
  output c0nm_b0m_wdata_3_;
  output c0nm_b0m_wdata_4_;
  output c0nm_b0m_wdata_5_;
  output c0nm_b0m_wdata_6_;
  output c0nm_b0m_wdata_7_;
  output c0nm_b0m_wdata_8_;
  output c0nm_b0m_wdata_9_;

  // moduleNum: x58
  // type: and2gate
  // conflicting modules: 
  // number of bit inputs: 11
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 1336/1336
  // type: INFERRED
  // marked bad? no
  // output word of size 10 : index:197 c0nm_b0m_wdata_11_ c0nm_b0m_wdata_8_ c0nm_b0m_wdata_9_ c0nm_b0m_wdata_7_
  // c0nm_b0m_wdata_6_ c0nm_b0m_wdata_5_ c0nm_b0m_wdata_4_ c0nm_b0m_wdata_3_ c0nm_b0m_wdata_2_ c0nm_b0m_wdata_10_
  // group: sel; nodes: [ c0nm_b0m_n1 ]

  AND2_X0P5M_A12TR c0nm_b0m_u13 (.A(flitin_0_10_), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_10_));
  AND2_X0P5M_A12TR c0nm_b0m_u12 (.A(flitin_0_11_), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_11_));
  AND2_X0P5M_A12TR c0nm_b0m_u11 (.A(flitin_0_2_), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_2_));
  AND2_X0P5M_A12TR c0nm_b0m_u10 (.A(flitin_0_3_), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_3_));
  AND2_X0P5M_A12TR c0nm_b0m_u9 (.A(flitin_0_4_), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_4_));
  AND2_X0P5M_A12TR c0nm_b0m_u8 (.A(flitin_0_5_), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_5_));
  AND2_X0P5M_A12TR c0nm_b0m_u7 (.A(flitin_0_6_), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_6_));
  AND2_X0P5M_A12TR c0nm_b0m_u6 (.A(flitin_0_7_), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_7_));
  AND2_X0P5M_A12TR c0nm_b0m_u5 (.A(flitin_0_8_), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_8_));
  AND2_X0P5M_A12TR c0nm_b0m_u4 (.A(flitin_0_9_), .B(c0nm_b0m_n1), .Y(c0nm_b0m_wdata_9_));
endmodule
module and2gate_mx59 
(
  c0nm_b0m_dqenablereg, 
  c0nm_b0m_rdata_10_, 
  c0nm_b0m_rdata_11_, 
  c0nm_b0m_rdata_2_, 
  c0nm_b0m_rdata_3_, 
  c0nm_b0m_rdata_4_, 
  c0nm_b0m_rdata_5_, 
  c0nm_b0m_rdata_6_, 
  c0nm_b0m_rdata_7_, 
  c0nm_b0m_rdata_8_, 
  c0nm_b0m_rdata_9_, 
  flitout_switch_0_10_,
  flitout_switch_0_11_,
  flitout_switch_0_2_,
  flitout_switch_0_3_,
  flitout_switch_0_4_,
  flitout_switch_0_5_,
  flitout_switch_0_6_,
  flitout_switch_0_7_,
  flitout_switch_0_8_,
  flitout_switch_0_9_
);
  input c0nm_b0m_dqenablereg;
  input c0nm_b0m_rdata_10_;
  input c0nm_b0m_rdata_11_;
  input c0nm_b0m_rdata_2_;
  input c0nm_b0m_rdata_3_;
  input c0nm_b0m_rdata_4_;
  input c0nm_b0m_rdata_5_;
  input c0nm_b0m_rdata_6_;
  input c0nm_b0m_rdata_7_;
  input c0nm_b0m_rdata_8_;
  input c0nm_b0m_rdata_9_;
  output flitout_switch_0_10_;
  output flitout_switch_0_11_;
  output flitout_switch_0_2_;
  output flitout_switch_0_3_;
  output flitout_switch_0_4_;
  output flitout_switch_0_5_;
  output flitout_switch_0_6_;
  output flitout_switch_0_7_;
  output flitout_switch_0_8_;
  output flitout_switch_0_9_;

  // moduleNum: x59
  // type: and2gate
  // conflicting modules: 
  // number of bit inputs: 11
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 1337/1337
  // type: INFERRED
  // marked bad? no
  // output word of size 10 : index:198 flitout_switch_0[11] flitout_switch_0[6] flitout_switch_0[5] flitout_switch_0[4]
  // flitout_switch_0[3] flitout_switch_0[2] flitout_switch_0[10] flitout_switch_0[9] flitout_switch_0[8] flitout_switch_0[7]
  // group: sel; nodes: [ c0nm_b0m_dqenablereg ]

  AND2_X0P5M_A12TR c0nm_b0m_u25 (.A(c0nm_b0m_rdata_10_), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0_10_));
  AND2_X0P5M_A12TR c0nm_b0m_u24 (.A(c0nm_b0m_rdata_11_), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0_11_));
  AND2_X0P5M_A12TR c0nm_b0m_u22 (.A(c0nm_b0m_rdata_2_), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0_2_));
  AND2_X0P5M_A12TR c0nm_b0m_u21 (.A(c0nm_b0m_rdata_3_), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0_3_));
  AND2_X0P5M_A12TR c0nm_b0m_u20 (.A(c0nm_b0m_rdata_4_), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0_4_));
  AND2_X0P5M_A12TR c0nm_b0m_u19 (.A(c0nm_b0m_rdata_5_), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0_5_));
  AND2_X0P5M_A12TR c0nm_b0m_u18 (.A(c0nm_b0m_rdata_6_), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0_6_));
  AND2_X0P5M_A12TR c0nm_b0m_u17 (.A(c0nm_b0m_rdata_7_), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0_7_));
  AND2_X0P5M_A12TR c0nm_b0m_u16 (.A(c0nm_b0m_rdata_8_), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0_8_));
  AND2_X0P5M_A12TR c0nm_b0m_u15 (.A(c0nm_b0m_rdata_9_), .B(c0nm_b0m_dqenablereg), .Y(flitout_switch_0_9_));
endmodule
module and2gate_mx60 
(
  c0nm_v0m_n5, 
  s0m_elig_1_, 
  swalloc_req_0_1_, 
  c0nm_v0m_n3,
  s0m_request0_1_
);
  input c0nm_v0m_n5;
  input s0m_elig_1_;
  input swalloc_req_0_1_;
  output c0nm_v0m_n3;
  output s0m_request0_1_;

  // moduleNum: x60
  // type: and2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1344/1346
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:200 s0m_request0[1] c0nm_v0m_n3 
  // group: sel; nodes: [ swalloc_req_0[1] ]

  AND2_X0P5M_A12TR c0nm_v0m_u5 (.A(swalloc_req_0_1_), .B(c0nm_v0m_n5), .Y(c0nm_v0m_n3));
  AND2_X0P5M_A12TR s0m_u10 (.A(s0m_elig_1_), .B(swalloc_req_0_1_), .Y(s0m_request0_1_));
endmodule
module and2gate_mx61 
(
  c0nm_v0m_n5, 
  s0m_elig_0_, 
  swalloc_req_0_0_, 
  c0nm_v0m_n7,
  s0m_request0_0_
);
  input c0nm_v0m_n5;
  input s0m_elig_0_;
  input swalloc_req_0_0_;
  output c0nm_v0m_n7;
  output s0m_request0_0_;

  // moduleNum: x61
  // type: and2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1347/1349
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:201 s0m_request0[0] c0nm_v0m_n7 
  // group: sel; nodes: [ swalloc_req_0[0] ]

  AND2_X0P5M_A12TR c0nm_v0m_u8 (.A(swalloc_req_0_0_), .B(c0nm_v0m_n5), .Y(c0nm_v0m_n7));
  AND2_X0P5M_A12TR s0m_u11 (.A(s0m_elig_0_), .B(swalloc_req_0_0_), .Y(s0m_request0_0_));
endmodule
module and2gate_mx62 
(
  c0sm_b0m_n2, 
  flitin_1_10_, 
  flitin_1_11_, 
  flitin_1_2_, 
  flitin_1_3_, 
  flitin_1_4_, 
  flitin_1_5_, 
  flitin_1_6_, 
  flitin_1_7_, 
  flitin_1_8_, 
  flitin_1_9_, 
  c0sm_b0m_wdata_10_,
  c0sm_b0m_wdata_11_,
  c0sm_b0m_wdata_2_,
  c0sm_b0m_wdata_3_,
  c0sm_b0m_wdata_4_,
  c0sm_b0m_wdata_5_,
  c0sm_b0m_wdata_6_,
  c0sm_b0m_wdata_7_,
  c0sm_b0m_wdata_8_,
  c0sm_b0m_wdata_9_
);
  input c0sm_b0m_n2;
  input flitin_1_10_;
  input flitin_1_11_;
  input flitin_1_2_;
  input flitin_1_3_;
  input flitin_1_4_;
  input flitin_1_5_;
  input flitin_1_6_;
  input flitin_1_7_;
  input flitin_1_8_;
  input flitin_1_9_;
  output c0sm_b0m_wdata_10_;
  output c0sm_b0m_wdata_11_;
  output c0sm_b0m_wdata_2_;
  output c0sm_b0m_wdata_3_;
  output c0sm_b0m_wdata_4_;
  output c0sm_b0m_wdata_5_;
  output c0sm_b0m_wdata_6_;
  output c0sm_b0m_wdata_7_;
  output c0sm_b0m_wdata_8_;
  output c0sm_b0m_wdata_9_;

  // moduleNum: x62
  // type: and2gate
  // conflicting modules: 
  // number of bit inputs: 11
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 1350/1350
  // type: INFERRED
  // marked bad? no
  // output word of size 10 : index:202 c0sm_b0m_wdata_10_ c0sm_b0m_wdata_9_ c0sm_b0m_wdata_8_ c0sm_b0m_wdata_7_
  // c0sm_b0m_wdata_6_ c0sm_b0m_wdata_5_ c0sm_b0m_wdata_4_ c0sm_b0m_wdata_3_ c0sm_b0m_wdata_11_ c0sm_b0m_wdata_2_
  // group: sel; nodes: [ c0sm_b0m_n2 ]

  AND2_X0P5M_A12TR c0sm_b0m_u13 (.A(flitin_1_10_), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_10_));
  AND2_X0P5M_A12TR c0sm_b0m_u12 (.A(flitin_1_11_), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_11_));
  AND2_X0P5M_A12TR c0sm_b0m_u11 (.A(flitin_1_2_), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_2_));
  AND2_X0P5M_A12TR c0sm_b0m_u10 (.A(flitin_1_3_), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_3_));
  AND2_X0P5M_A12TR c0sm_b0m_u9 (.A(flitin_1_4_), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_4_));
  AND2_X0P5M_A12TR c0sm_b0m_u8 (.A(flitin_1_5_), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_5_));
  AND2_X0P5M_A12TR c0sm_b0m_u7 (.A(flitin_1_6_), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_6_));
  AND2_X0P5M_A12TR c0sm_b0m_u6 (.A(flitin_1_7_), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_7_));
  AND2_X0P5M_A12TR c0sm_b0m_u5 (.A(flitin_1_8_), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_8_));
  AND2_X0P5M_A12TR c0sm_b0m_u4 (.A(flitin_1_9_), .B(c0sm_b0m_n2), .Y(c0sm_b0m_wdata_9_));
endmodule
module and2gate_mx63 
(
  c0sm_b0m_dqenablereg, 
  c0sm_b0m_rdata_10_, 
  c0sm_b0m_rdata_11_, 
  c0sm_b0m_rdata_2_, 
  c0sm_b0m_rdata_3_, 
  c0sm_b0m_rdata_4_, 
  c0sm_b0m_rdata_5_, 
  c0sm_b0m_rdata_6_, 
  c0sm_b0m_rdata_7_, 
  c0sm_b0m_rdata_8_, 
  c0sm_b0m_rdata_9_, 
  flitout_switch_1_10_,
  flitout_switch_1_11_,
  flitout_switch_1_2_,
  flitout_switch_1_3_,
  flitout_switch_1_4_,
  flitout_switch_1_5_,
  flitout_switch_1_6_,
  flitout_switch_1_7_,
  flitout_switch_1_8_,
  flitout_switch_1_9_
);
  input c0sm_b0m_dqenablereg;
  input c0sm_b0m_rdata_10_;
  input c0sm_b0m_rdata_11_;
  input c0sm_b0m_rdata_2_;
  input c0sm_b0m_rdata_3_;
  input c0sm_b0m_rdata_4_;
  input c0sm_b0m_rdata_5_;
  input c0sm_b0m_rdata_6_;
  input c0sm_b0m_rdata_7_;
  input c0sm_b0m_rdata_8_;
  input c0sm_b0m_rdata_9_;
  output flitout_switch_1_10_;
  output flitout_switch_1_11_;
  output flitout_switch_1_2_;
  output flitout_switch_1_3_;
  output flitout_switch_1_4_;
  output flitout_switch_1_5_;
  output flitout_switch_1_6_;
  output flitout_switch_1_7_;
  output flitout_switch_1_8_;
  output flitout_switch_1_9_;

  // moduleNum: x63
  // type: and2gate
  // conflicting modules: 
  // number of bit inputs: 11
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 10
  // number of non-inferred gates: 0
  // ILP vars: 1351/1351
  // type: INFERRED
  // marked bad? no
  // output word of size 10 : index:203 flitout_switch_1[5] flitout_switch_1[9] flitout_switch_1[8] flitout_switch_1[7]
  // flitout_switch_1[6] flitout_switch_1[4] flitout_switch_1[3] flitout_switch_1[2] flitout_switch_1[11]
  // flitout_switch_1[10]
  // group: sel; nodes: [ c0sm_b0m_dqenablereg ]

  AND2_X0P5M_A12TR c0sm_b0m_u25 (.A(c0sm_b0m_rdata_10_), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1_10_));
  AND2_X0P5M_A12TR c0sm_b0m_u24 (.A(c0sm_b0m_rdata_11_), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1_11_));
  AND2_X0P5M_A12TR c0sm_b0m_u22 (.A(c0sm_b0m_rdata_2_), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1_2_));
  AND2_X0P5M_A12TR c0sm_b0m_u21 (.A(c0sm_b0m_rdata_3_), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1_3_));
  AND2_X0P5M_A12TR c0sm_b0m_u20 (.A(c0sm_b0m_rdata_4_), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1_4_));
  AND2_X0P5M_A12TR c0sm_b0m_u19 (.A(c0sm_b0m_rdata_5_), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1_5_));
  AND2_X0P5M_A12TR c0sm_b0m_u18 (.A(c0sm_b0m_rdata_6_), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1_6_));
  AND2_X0P5M_A12TR c0sm_b0m_u17 (.A(c0sm_b0m_rdata_7_), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1_7_));
  AND2_X0P5M_A12TR c0sm_b0m_u16 (.A(c0sm_b0m_rdata_8_), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1_8_));
  AND2_X0P5M_A12TR c0sm_b0m_u15 (.A(c0sm_b0m_rdata_9_), .B(c0sm_b0m_dqenablereg), .Y(flitout_switch_1_9_));
endmodule
module and2gate_mx64 
(
  c0sm_v0m_n5, 
  s0m_elig_1_, 
  swalloc_req_1_1_, 
  c0sm_v0m_n3,
  s0m_request1_1_
);
  input c0sm_v0m_n5;
  input s0m_elig_1_;
  input swalloc_req_1_1_;
  output c0sm_v0m_n3;
  output s0m_request1_1_;

  // moduleNum: x64
  // type: and2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1358/1360
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:206 s0m_request1[1] c0sm_v0m_n3 
  // group: sel; nodes: [ swalloc_req_1[1] ]

  AND2_X0P5M_A12TR c0sm_v0m_u5 (.A(swalloc_req_1_1_), .B(c0sm_v0m_n5), .Y(c0sm_v0m_n3));
  AND2_X0P5M_A12TR s0m_u8 (.A(s0m_elig_1_), .B(swalloc_req_1_1_), .Y(s0m_request1_1_));
endmodule
module and2gate_mx65 
(
  c0sm_v0m_n5, 
  s0m_elig_0_, 
  swalloc_req_1_0_, 
  c0sm_v0m_n7,
  s0m_request1_0_
);
  input c0sm_v0m_n5;
  input s0m_elig_0_;
  input swalloc_req_1_0_;
  output c0sm_v0m_n7;
  output s0m_request1_0_;

  // moduleNum: x65
  // type: and2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1361/1363
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:207 s0m_request1[0] c0sm_v0m_n7 
  // group: sel; nodes: [ swalloc_req_1[0] ]

  AND2_X0P5M_A12TR c0sm_v0m_u8 (.A(swalloc_req_1_0_), .B(c0sm_v0m_n5), .Y(c0sm_v0m_n7));
  AND2_X0P5M_A12TR s0m_u9 (.A(s0m_elig_0_), .B(swalloc_req_1_0_), .Y(s0m_request1_0_));
endmodule
module or2gate_mx66 
(
  c0nm_r0m_n9, 
  c0sm_r0m_n9, 
  currx_0_, 
  c0nm_r0m_n15,
  c0sm_r0m_n15
);
  input c0nm_r0m_n9;
  input c0sm_r0m_n9;
  input currx_0_;
  output c0nm_r0m_n15;
  output c0sm_r0m_n15;

  // moduleNum: x66
  // type: or2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1370/1370
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:210 c0nm_r0m_n15 c0sm_r0m_n15 
  // group: sel; nodes: [ currx[0] ]

  OR2_X0P5M_A12TR c0nm_r0m_u18 (.A(currx_0_), .B(c0nm_r0m_n9), .Y(c0nm_r0m_n15));
  OR2_X0P5M_A12TR c0sm_r0m_u18 (.A(currx_0_), .B(c0sm_r0m_n9), .Y(c0sm_r0m_n15));
endmodule
module or2gate_mx67 
(
  c0nm_b0m_n1, 
  c0nm_b0m_v0m_n8, 
  c0nm_b0m_v0m_n93, 
  c0nm_b0m_v0m_n94, 
  c0nm_b0m_v0m_n95, 
  c0nm_headflit_0_, 
  c0nm_headflit_1_, 
  c0sm_b0m_n2, 
  c0sm_b0m_v0m_n8, 
  c0sm_b0m_v0m_n93, 
  c0sm_b0m_v0m_n94, 
  c0sm_b0m_v0m_n95, 
  c0sm_headflit_0_, 
  c0sm_headflit_1_, 
  colsel0_0_, 
  colsel0_1_, 
  colsel1_0_, 
  colsel1_1_, 
  reset, 
  tailout_0, 
  tailout_1, 
  c0nm_b0m_v0m_n1,
  c0nm_b0m_v0m_n102,
  c0nm_b0m_v0m_n129,
  c0nm_b0m_v0m_n2,
  c0nm_b0m_v0m_n262,
  c0nm_b0m_v0m_n263,
  c0nm_b0m_v0m_n81,
  c0nm_v0m_n1,
  c0sm_b0m_v0m_n1,
  c0sm_b0m_v0m_n102,
  c0sm_b0m_v0m_n129,
  c0sm_b0m_v0m_n2,
  c0sm_b0m_v0m_n262,
  c0sm_b0m_v0m_n263,
  c0sm_b0m_v0m_n81,
  c0sm_v0m_n1,
  x0m_n3,
  x0m_n4,
  x0m_n5,
  x0m_n6
);
  input c0nm_b0m_n1;
  input c0nm_b0m_v0m_n8;
  input c0nm_b0m_v0m_n93;
  input c0nm_b0m_v0m_n94;
  input c0nm_b0m_v0m_n95;
  input c0nm_headflit_0_;
  input c0nm_headflit_1_;
  input c0sm_b0m_n2;
  input c0sm_b0m_v0m_n8;
  input c0sm_b0m_v0m_n93;
  input c0sm_b0m_v0m_n94;
  input c0sm_b0m_v0m_n95;
  input c0sm_headflit_0_;
  input c0sm_headflit_1_;
  input colsel0_0_;
  input colsel0_1_;
  input colsel1_0_;
  input colsel1_1_;
  input reset;
  input tailout_0;
  input tailout_1;
  output c0nm_b0m_v0m_n1;
  output c0nm_b0m_v0m_n102;
  output c0nm_b0m_v0m_n129;
  output c0nm_b0m_v0m_n2;
  output c0nm_b0m_v0m_n262;
  output c0nm_b0m_v0m_n263;
  output c0nm_b0m_v0m_n81;
  output c0nm_v0m_n1;
  output c0sm_b0m_v0m_n1;
  output c0sm_b0m_v0m_n102;
  output c0sm_b0m_v0m_n129;
  output c0sm_b0m_v0m_n2;
  output c0sm_b0m_v0m_n262;
  output c0sm_b0m_v0m_n263;
  output c0sm_b0m_v0m_n81;
  output c0sm_v0m_n1;
  output x0m_n3;
  output x0m_n4;
  output x0m_n5;
  output x0m_n6;
  wire c0nm_b0m_v0m_n108;
  wire c0nm_b0m_v0m_n264;
  wire c0nm_b0m_v0m_n4;
  wire c0nm_b0m_v0m_n77;
  wire c0nm_b0m_v0m_n99;
  wire c0nm_v0m_n8;
  wire c0sm_b0m_v0m_n108;
  wire c0sm_b0m_v0m_n264;
  wire c0sm_b0m_v0m_n77;
  wire c0sm_b0m_v0m_n99;
  wire c0sm_v0m_n8;

  // moduleNum: x67
  // type: or2gate
  // conflicting modules: 
  // number of bit inputs: 21
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 31
  // number of non-inferred gates: 0
  // ILP vars: 1371/1371
  // type: INFERRED
  // marked bad? no
  // output word of size 20 : index:211 x0m_n3 x0m_n4 x0m_n5 x0m_n6 c0nm_v0m_n1 c0sm_v0m_n1 c0sm_b0m_v0m_n1 c0nm_b0m_v0m_n1
  // c0sm_b0m_v0m_n81 c0sm_b0m_v0m_n2 c0sm_b0m_v0m_n129 c0sm_b0m_v0m_n102 c0nm_b0m_v0m_n2 c0nm_b0m_v0m_n81 c0nm_b0m_v0m_n102
  // c0nm_b0m_v0m_n129 c0sm_b0m_v0m_n262 c0nm_b0m_v0m_n262 c0nm_b0m_v0m_n263 c0sm_b0m_v0m_n263
  // group: sel; nodes: [ reset ]

  INV_X0P5B_A12TR c0nm_b0m_v0m_u262 (.A(c0nm_headflit_1_), .Y(c0nm_b0m_v0m_n264));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u261 (.A(reset), .Y(c0nm_b0m_v0m_n4));
  NAND2_X0P5A_A12TR c0nm_b0m_v0m_u197 (.A(c0nm_b0m_v0m_n264), .B(c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n263));
  NAND2B_X0P5M_A12TR c0nm_b0m_v0m_u195 (.AN(c0nm_headflit_0_), .B(c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n262));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u179 (.A(c0nm_b0m_v0m_n94), .Y(c0nm_b0m_v0m_n108));
  NAND2_X0P5A_A12TR c0nm_b0m_v0m_u178 (.A(c0nm_b0m_v0m_n108), .B(c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n129));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u83 (.A(c0nm_b0m_v0m_n93), .Y(c0nm_b0m_v0m_n99));
  NAND2_X0P5A_A12TR c0nm_b0m_v0m_u82 (.A(c0nm_b0m_v0m_n99), .B(c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n102));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u64 (.A(c0nm_b0m_v0m_n95), .Y(c0nm_b0m_v0m_n77));
  NAND2_X0P5A_A12TR c0nm_b0m_v0m_u63 (.A(c0nm_b0m_v0m_n77), .B(c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n81));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u7 (.A(c0nm_b0m_v0m_n8), .Y(c0nm_b0m_v0m_n1));
  NAND2_X0P5A_A12TR c0nm_b0m_v0m_u4 (.A(c0nm_b0m_v0m_n1), .B(c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n2));
  NOR2_X0P5A_A12TR c0nm_v0m_u38 (.A(reset), .B(tailout_0), .Y(c0nm_v0m_n8));
  INV_X0P5B_A12TR c0nm_v0m_u9 (.A(c0nm_v0m_n8), .Y(c0nm_v0m_n1));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u262 (.A(c0sm_headflit_1_), .Y(c0sm_b0m_v0m_n264));
  NAND2_X0P5A_A12TR c0sm_b0m_v0m_u197 (.A(c0sm_b0m_v0m_n264), .B(c0nm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n263));
  NAND2B_X0P5M_A12TR c0sm_b0m_v0m_u195 (.AN(c0sm_headflit_0_), .B(c0nm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n262));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u179 (.A(c0sm_b0m_v0m_n94), .Y(c0sm_b0m_v0m_n108));
  NAND2_X0P5A_A12TR c0sm_b0m_v0m_u178 (.A(c0sm_b0m_v0m_n108), .B(c0nm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n129));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u83 (.A(c0sm_b0m_v0m_n93), .Y(c0sm_b0m_v0m_n99));
  NAND2_X0P5A_A12TR c0sm_b0m_v0m_u82 (.A(c0sm_b0m_v0m_n99), .B(c0nm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n102));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u64 (.A(c0sm_b0m_v0m_n95), .Y(c0sm_b0m_v0m_n77));
  NAND2_X0P5A_A12TR c0sm_b0m_v0m_u63 (.A(c0sm_b0m_v0m_n77), .B(c0nm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n81));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u7 (.A(c0sm_b0m_v0m_n8), .Y(c0sm_b0m_v0m_n1));
  NAND2_X0P5A_A12TR c0sm_b0m_v0m_u4 (.A(c0sm_b0m_v0m_n1), .B(c0nm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n2));
  NOR2_X0P5A_A12TR c0sm_v0m_u38 (.A(reset), .B(tailout_1), .Y(c0sm_v0m_n8));
  INV_X0P5B_A12TR c0sm_v0m_u9 (.A(c0sm_v0m_n8), .Y(c0sm_v0m_n1));
  OR2_X0P5M_A12TR x0m_u8 (.A(colsel0_0_), .B(reset), .Y(x0m_n3));
  OR2_X0P5M_A12TR x0m_u7 (.A(colsel0_1_), .B(reset), .Y(x0m_n4));
  OR2_X0P5M_A12TR x0m_u6 (.A(colsel1_0_), .B(reset), .Y(x0m_n5));
  OR2_X0P5M_A12TR x0m_u5 (.A(colsel1_1_), .B(reset), .Y(x0m_n6));
endmodule
module or2gate_mx68 
(
  c0nm_b0m_n1, 
  c0nm_b0m_v0m_n28, 
  c0nm_b0m_v0m_n93, 
  c0nm_b0m_v0m_n116,
  c0nm_b0m_v0m_n135
);
  input c0nm_b0m_n1;
  input c0nm_b0m_v0m_n28;
  input c0nm_b0m_v0m_n93;
  output c0nm_b0m_v0m_n116;
  output c0nm_b0m_v0m_n135;
  wire c0nm_b0m_v0m_n119;
  wire c0nm_b0m_v0m_n128;

  // moduleNum: x68
  // type: or2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 4
  // number of non-inferred gates: 0
  // ILP vars: 1372/1375
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:246 c0nm_b0m_v0m_n135 c0nm_b0m_v0m_n116 
  // group: sel; nodes: [ c0nm_b0m_n1 ]

  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u191 (.A(c0nm_b0m_v0m_n93), .B(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n119));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u190 (.A(c0nm_b0m_v0m_n119), .Y(c0nm_b0m_v0m_n135));
  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u182 (.A(c0nm_b0m_v0m_n28), .B(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n128));
  INV_X0P5B_A12TR c0nm_b0m_v0m_u98 (.A(c0nm_b0m_v0m_n128), .Y(c0nm_b0m_v0m_n116));
endmodule
module or2gate_mx69 
(
  c0sm_b0m_n2, 
  c0sm_b0m_v0m_n28, 
  c0sm_b0m_v0m_n93, 
  c0sm_b0m_v0m_n116,
  c0sm_b0m_v0m_n135
);
  input c0sm_b0m_n2;
  input c0sm_b0m_v0m_n28;
  input c0sm_b0m_v0m_n93;
  output c0sm_b0m_v0m_n116;
  output c0sm_b0m_v0m_n135;
  wire c0sm_b0m_v0m_n119;
  wire c0sm_b0m_v0m_n128;

  // moduleNum: x69
  // type: or2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 4
  // number of non-inferred gates: 0
  // ILP vars: 1379/1382
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:247 c0sm_b0m_v0m_n135 c0sm_b0m_v0m_n116 
  // group: sel; nodes: [ c0sm_b0m_n2 ]

  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u191 (.A(c0sm_b0m_v0m_n93), .B(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n119));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u190 (.A(c0sm_b0m_v0m_n119), .Y(c0sm_b0m_v0m_n135));
  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u182 (.A(c0sm_b0m_v0m_n28), .B(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n128));
  INV_X0P5B_A12TR c0sm_b0m_v0m_u98 (.A(c0sm_b0m_v0m_n128), .Y(c0sm_b0m_v0m_n116));
endmodule
module or2gate_mx70 
(
  x0m_bx0m_m1m_int01, 
  x0m_bx1m_m1m_int01, 
  x0m_colsel1reg_1_, 
  flitout_1_0_,
  flitout_1_1_
);
  input x0m_bx0m_m1m_int01;
  input x0m_bx1m_m1m_int01;
  input x0m_colsel1reg_1_;
  output flitout_1_0_;
  output flitout_1_1_;
  wire x0m__logic1_;

  // moduleNum: x70
  // type: or2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 3
  // number of non-inferred gates: 0
  // ILP vars: 1389/1391
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:217 flitout_1[1] flitout_1[0] 
  // group: sel; nodes: [ x0m_colsel1reg_1_ ]

  TIEHI_X1M_A12TR x0m_u4 (.Y(x0m__logic1_));
  MXT2_X0P5M_A12TR x0m_bx0m_m1m_m4m_u1 (.A(x0m_bx0m_m1m_int01), .B(x0m__logic1_), .S0(x0m_colsel1reg_1_), .Y(flitout_1_0_));
  MXT2_X0P5M_A12TR x0m_bx1m_m1m_m4m_u1 (.A(x0m_bx1m_m1m_int01), .B(x0m__logic1_), .S0(x0m_colsel1reg_1_), .Y(flitout_1_1_));
endmodule
module nand2gate_mx71 
(
  flitin_0_0_, 
  flitin_0_1_, 
  c0nm_b0m_n1,
  c0nm_n2
);
  input flitin_0_0_;
  input flitin_0_1_;
  output c0nm_b0m_n1;
  output c0nm_n2;

  // moduleNum: x71
  // type: nand2gate
  // conflicting modules: 
  // number of bit inputs: 2
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1395/1397
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:-1 c0nm_n2 c0nm_b0m_n1 
  // group: sel; nodes: [ flitin_0[0] ]

  NAND2_X0P5A_A12TR c0nm_u3 (.A(flitin_0_1_), .B(flitin_0_0_), .Y(c0nm_n2));
  NAND2_X0P5A_A12TR c0nm_b0m_u14 (.A(flitin_0_1_), .B(flitin_0_0_), .Y(c0nm_b0m_n1));
endmodule
module nand2gate_mx72 
(
  flitin_1_0_, 
  flitin_1_1_, 
  c0sm_b0m_n2,
  c0sm_n3
);
  input flitin_1_0_;
  input flitin_1_1_;
  output c0sm_b0m_n2;
  output c0sm_n3;

  // moduleNum: x72
  // type: nand2gate
  // conflicting modules: 
  // number of bit inputs: 2
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1401/1403
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:-1 c0sm_n3 c0sm_b0m_n2 
  // group: sel; nodes: [ flitin_1[0] ]

  NAND2_X0P5A_A12TR c0sm_u3 (.A(flitin_1_1_), .B(flitin_1_0_), .Y(c0sm_n3));
  NAND2_X0P5A_A12TR c0sm_b0m_u14 (.A(flitin_1_1_), .B(flitin_1_0_), .Y(c0sm_b0m_n2));
endmodule
module nand2gate_mx73 
(
  c0nm_b0m_v0m_n26, 
  c0nm_b0m_v0m_n4, 
  c0sm_b0m_v0m_n26, 
  s0m_o0nm_n24, 
  s0m_o0sm_n24, 
  c0nm_b0m_v0m_n20,
  c0sm_b0m_v0m_n20,
  s0m_o0nm_n36,
  s0m_o0sm_n36
);
  input c0nm_b0m_v0m_n26;
  input c0nm_b0m_v0m_n4;
  input c0sm_b0m_v0m_n26;
  input s0m_o0nm_n24;
  input s0m_o0sm_n24;
  output c0nm_b0m_v0m_n20;
  output c0sm_b0m_v0m_n20;
  output s0m_o0nm_n36;
  output s0m_o0sm_n36;

  // moduleNum: x73
  // type: nand2gate
  // conflicting modules: 
  // number of bit inputs: 5
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 4
  // number of non-inferred gates: 0
  // ILP vars: 1404/1418
  // type: INFERRED
  // marked bad? no
  // output word of size 4 : index:248 c0sm_b0m_v0m_n20 c0nm_b0m_v0m_n20 s0m_o0nm_n36 s0m_o0sm_n36 
  // group: sel; nodes: [ c0nm_b0m_v0m_n4 ]

  NAND2_X0P5A_A12TR c0nm_b0m_v0m_u31 (.A(c0nm_b0m_v0m_n26), .B(c0nm_b0m_v0m_n4), .Y(c0nm_b0m_v0m_n20));
  NAND2_X0P5A_A12TR c0sm_b0m_v0m_u31 (.A(c0sm_b0m_v0m_n26), .B(c0nm_b0m_v0m_n4), .Y(c0sm_b0m_v0m_n20));
  NAND2_X0P5A_A12TR s0m_o0nm_u23 (.A(s0m_o0nm_n24), .B(c0nm_b0m_v0m_n4), .Y(s0m_o0nm_n36));
  NAND2_X0P5A_A12TR s0m_o0sm_u23 (.A(s0m_o0sm_n24), .B(c0nm_b0m_v0m_n4), .Y(s0m_o0sm_n36));
endmodule
module nand2gate_mx74 
(
  s0m_state_invc0_1_, 
  s0m_state_invc1_1_, 
  tailout_1, 
  s0m_n1,
  s0m_n3
);
  input s0m_state_invc0_1_;
  input s0m_state_invc1_1_;
  input tailout_1;
  output s0m_n1;
  output s0m_n3;

  // moduleNum: x74
  // type: nand2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1419/1421
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:221 s0m_n3 s0m_n1 
  // group: sel; nodes: [ tailout_1 ]

  NAND2_X0P5A_A12TR s0m_u7 (.A(s0m_state_invc0_1_), .B(tailout_1), .Y(s0m_n3));
  NAND2_X0P5A_A12TR s0m_u4 (.A(tailout_1), .B(s0m_state_invc1_1_), .Y(s0m_n1));
endmodule
module nand2gate_mx75 
(
  debitout_1, 
  s0m_state_invc0_1_, 
  s0m_state_invc1_1_, 
  s0m_n20,
  s0m_n26
);
  input debitout_1;
  input s0m_state_invc0_1_;
  input s0m_state_invc1_1_;
  output s0m_n20;
  output s0m_n26;

  // moduleNum: x75
  // type: nand2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1422/1424
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:222 s0m_n26 s0m_n20 
  // group: sel; nodes: [ debitout_1 ]

  NAND2_X0P5A_A12TR s0m_u38 (.A(debitout_1), .B(s0m_state_invc0_1_), .Y(s0m_n26));
  NAND2_X0P5A_A12TR s0m_u35 (.A(debitout_1), .B(s0m_state_invc1_1_), .Y(s0m_n20));
endmodule
module nand2gate_mx76 
(
  s0m_n16, 
  s0m_outb0_1_, 
  s0m_outb1_1_, 
  s0m_n14,
  s0m_n18
);
  input s0m_n16;
  input s0m_outb0_1_;
  input s0m_outb1_1_;
  output s0m_n14;
  output s0m_n18;

  // moduleNum: x76
  // type: nand2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1425/1425
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:223 s0m_n18 s0m_n14 
  // group: sel; nodes: [ s0m_n16 ]

  NAND2_X0P5A_A12TR s0m_u31 (.A(s0m_outb1_1_), .B(s0m_n16), .Y(s0m_n18));
  NAND2_X0P5A_A12TR s0m_u26 (.A(s0m_outb0_1_), .B(s0m_n16), .Y(s0m_n14));
endmodule
module nand2gate_mx77 
(
  s0m_n9, 
  s0m_outb0_0_, 
  s0m_outb1_0_, 
  s0m_n11,
  s0m_n7
);
  input s0m_n9;
  input s0m_outb0_0_;
  input s0m_outb1_0_;
  output s0m_n11;
  output s0m_n7;

  // moduleNum: x77
  // type: nand2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1426/1426
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:224 s0m_n11 s0m_n7 
  // group: sel; nodes: [ s0m_n9 ]

  NAND2_X0P5A_A12TR s0m_u22 (.A(s0m_outb1_0_), .B(s0m_n9), .Y(s0m_n11));
  NAND2_X0P5A_A12TR s0m_u17 (.A(s0m_outb0_0_), .B(s0m_n9), .Y(s0m_n7));
endmodule
module nor2gate_mx78 
(
  c0nm_b0m_n1, 
  c0nm_v0m_n10, 
  c0nm_v0m_n19, 
  c0nm_v0m_n27, 
  c0sm_b0m_n2, 
  c0sm_v0m_n10, 
  c0sm_v0m_n19, 
  c0sm_v0m_n27, 
  debitout_0, 
  debitout_1, 
  reset, 
  s0m_m0m_n2, 
  s0m_m1m_n2, 
  s0m_o0nm_n13, 
  s0m_o0sm_n13, 
  s0m_tail_outvc0, 
  s0m_tail_outvc1, 
  tailout_0, 
  tailout_1, 
  c0nm_b0m_v0m_n10,
  c0nm_b0m_v0m_n11,
  c0nm_b0m_v0m_n8,
  c0nm_v0m_n61,
  c0nm_v0m_n62,
  c0nm_v0m_n64,
  c0sm_b0m_v0m_n10,
  c0sm_b0m_v0m_n11,
  c0sm_b0m_v0m_n8,
  c0sm_v0m_n61,
  c0sm_v0m_n62,
  c0sm_v0m_n64,
  creditout_0,
  creditout_1,
  s0m_m0m_n10,
  s0m_m1m_n10,
  s0m_n16,
  s0m_n9,
  s0m_o0nm_n3,
  s0m_o0nm_n38,
  s0m_o0sm_n3,
  s0m_o0sm_n38
);
  input c0nm_b0m_n1;
  input c0nm_v0m_n10;
  input c0nm_v0m_n19;
  input c0nm_v0m_n27;
  input c0sm_b0m_n2;
  input c0sm_v0m_n10;
  input c0sm_v0m_n19;
  input c0sm_v0m_n27;
  input debitout_0;
  input debitout_1;
  input reset;
  input s0m_m0m_n2;
  input s0m_m1m_n2;
  input s0m_o0nm_n13;
  input s0m_o0sm_n13;
  input s0m_tail_outvc0;
  input s0m_tail_outvc1;
  input tailout_0;
  input tailout_1;
  output c0nm_b0m_v0m_n10;
  output c0nm_b0m_v0m_n11;
  output c0nm_b0m_v0m_n8;
  output c0nm_v0m_n61;
  output c0nm_v0m_n62;
  output c0nm_v0m_n64;
  output c0sm_b0m_v0m_n10;
  output c0sm_b0m_v0m_n11;
  output c0sm_b0m_v0m_n8;
  output c0sm_v0m_n61;
  output c0sm_v0m_n62;
  output c0sm_v0m_n64;
  output creditout_0;
  output creditout_1;
  output s0m_m0m_n10;
  output s0m_m1m_n10;
  output s0m_n16;
  output s0m_n9;
  output s0m_o0nm_n3;
  output s0m_o0nm_n38;
  output s0m_o0sm_n3;
  output s0m_o0sm_n38;

  // moduleNum: x78
  // type: nor2gate
  // conflicting modules: 
  // number of bit inputs: 19
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 22
  // number of non-inferred gates: 0
  // ILP vars: 1433/1463
  // type: INFERRED
  // marked bad? no
  // output word of size 26 : index:249 s0m_n9 s0m_n16 c0nm_b0m_v0m_n8 c0sm_b0m_v0m_n8 s0m_o0nm_n3 s0m_o0sm_n3 s0m_m0m_n10
  // s0m_m0m_n10 c0nm_b0m_v0m_n11 c0sm_b0m_v0m_n11 s0m_m1m_n10 s0m_m1m_n10 creditout_0 creditout_1 c0sm_b0m_v0m_n10
  // c0sm_b0m_v0m_n10 c0nm_b0m_v0m_n10 c0nm_b0m_v0m_n10 c0sm_v0m_n64 c0nm_v0m_n64 c0sm_v0m_n61 c0nm_v0m_n61 c0sm_v0m_n62
  // c0nm_v0m_n62 s0m_o0nm_n38 s0m_o0sm_n38
  // group: sel; nodes: [ reset ]

  NOR2B_X0P5M_A12TR c0nm_u5 (.AN(debitout_0), .B(reset), .Y(creditout_0));
  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u209 (.A(debitout_0), .B(reset), .Y(c0nm_b0m_v0m_n11));
  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u208 (.A(c0nm_b0m_v0m_n11), .B(reset), .Y(c0nm_b0m_v0m_n10));
  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u10 (.A(reset), .B(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n8));
  NOR2_X0P5A_A12TR c0nm_v0m_u23 (.A(reset), .B(c0nm_v0m_n27), .Y(c0nm_v0m_n61));
  NOR2_X0P5A_A12TR c0nm_v0m_u17 (.A(reset), .B(c0nm_v0m_n19), .Y(c0nm_v0m_n62));
  NOR2_X0P5A_A12TR c0nm_v0m_u11 (.A(reset), .B(c0nm_v0m_n10), .Y(c0nm_v0m_n64));
  NOR2B_X0P5M_A12TR c0sm_u5 (.AN(debitout_1), .B(reset), .Y(creditout_1));
  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u209 (.A(debitout_1), .B(reset), .Y(c0sm_b0m_v0m_n11));
  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u208 (.A(c0sm_b0m_v0m_n11), .B(reset), .Y(c0sm_b0m_v0m_n10));
  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u10 (.A(reset), .B(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n8));
  NOR2_X0P5A_A12TR c0sm_v0m_u23 (.A(reset), .B(c0sm_v0m_n27), .Y(c0sm_v0m_n61));
  NOR2_X0P5A_A12TR c0sm_v0m_u17 (.A(reset), .B(c0sm_v0m_n19), .Y(c0sm_v0m_n62));
  NOR2_X0P5A_A12TR c0sm_v0m_u11 (.A(reset), .B(c0sm_v0m_n10), .Y(c0sm_v0m_n64));
  NOR2_X0P5A_A12TR s0m_u32 (.A(reset), .B(tailout_1), .Y(s0m_n16));
  NOR2_X0P5A_A12TR s0m_u23 (.A(reset), .B(tailout_0), .Y(s0m_n9));
  NOR2_X0P5A_A12TR s0m_m0m_u4 (.A(reset), .B(s0m_m0m_n2), .Y(s0m_m0m_n10));
  NOR2_X0P5A_A12TR s0m_m1m_u4 (.A(reset), .B(s0m_m1m_n2), .Y(s0m_m1m_n10));
  NOR2_X0P5A_A12TR s0m_o0nm_u35 (.A(s0m_tail_outvc0), .B(reset), .Y(s0m_o0nm_n3));
  NOR2_X0P5A_A12TR s0m_o0nm_u14 (.A(reset), .B(s0m_o0nm_n13), .Y(s0m_o0nm_n38));
  NOR2_X0P5A_A12TR s0m_o0sm_u35 (.A(s0m_tail_outvc1), .B(reset), .Y(s0m_o0sm_n3));
  NOR2_X0P5A_A12TR s0m_o0sm_u14 (.A(reset), .B(s0m_o0sm_n13), .Y(s0m_o0sm_n38));
endmodule
module nor2gate_mx79 
(
  c0nm_b0m_n1, 
  c0nm_b0m_v0m_n94, 
  c0nm_b0m_v0m_n95, 
  c0nm_b0m_v0m_n120,
  c0nm_b0m_v0m_n121
);
  input c0nm_b0m_n1;
  input c0nm_b0m_v0m_n94;
  input c0nm_b0m_v0m_n95;
  output c0nm_b0m_v0m_n120;
  output c0nm_b0m_v0m_n121;

  // moduleNum: x79
  // type: nor2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1464/1469
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:250 c0nm_b0m_v0m_n120 c0nm_b0m_v0m_n121 
  // group: sel; nodes: [ c0nm_b0m_n1 ]

  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u187 (.A(c0nm_b0m_v0m_n94), .B(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n121));
  NOR2_X0P5A_A12TR c0nm_b0m_v0m_u185 (.A(c0nm_b0m_v0m_n95), .B(c0nm_b0m_n1), .Y(c0nm_b0m_v0m_n120));
endmodule
module nor2gate_mx80 
(
  c0nm_n2, 
  c0nm_v0m_n9, 
  reset, 
  c0nm_b0m_n9,
  c0nm_v0m_n13
);
  input c0nm_n2;
  input c0nm_v0m_n9;
  input reset;
  output c0nm_b0m_n9;
  output c0nm_v0m_n13;
  wire debitout_0;

  // moduleNum: x80
  // type: nor2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 3
  // number of non-inferred gates: 0
  // ILP vars: 1473/1477
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:251 c0nm_v0m_n13 c0nm_b0m_n9 
  // group: sel; nodes: [ c0nm_v0m_n9 ]

  NOR2B_X0P5M_A12TR c0nm_b0m_u27 (.AN(debitout_0), .B(reset), .Y(c0nm_b0m_n9));
  NOR2_X0P5A_A12TR c0nm_v0m_u30 (.A(c0nm_v0m_n9), .B(c0nm_n2), .Y(c0nm_v0m_n13));
  INV_X0P5B_A12TR c0nm_v0m_u10 (.A(c0nm_v0m_n9), .Y(debitout_0));
endmodule
module nor2gate_mx81 
(
  c0nm_v0m_n1, 
  c0nm_v0m_n2, 
  c0nm_v0m_n6, 
  c0nm_v0m_n30,
  c0nm_v0m_n31
);
  input c0nm_v0m_n1;
  input c0nm_v0m_n2;
  input c0nm_v0m_n6;
  output c0nm_v0m_n30;
  output c0nm_v0m_n31;

  // moduleNum: x81
  // type: nor2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1482/1482
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:231 c0nm_v0m_n31 c0nm_v0m_n30 
  // group: sel; nodes: [ c0nm_v0m_n1 ]

  NOR2_X0P5A_A12TR c0nm_v0m_u6 (.A(c0nm_v0m_n1), .B(c0nm_v0m_n6), .Y(c0nm_v0m_n30));
  NOR2_X0P5A_A12TR c0nm_v0m_u3 (.A(c0nm_v0m_n1), .B(c0nm_v0m_n2), .Y(c0nm_v0m_n31));
endmodule
module nor2gate_mx82 
(
  c0sm_b0m_n2, 
  c0sm_b0m_v0m_n94, 
  c0sm_b0m_v0m_n95, 
  c0sm_b0m_v0m_n120,
  c0sm_b0m_v0m_n121
);
  input c0sm_b0m_n2;
  input c0sm_b0m_v0m_n94;
  input c0sm_b0m_v0m_n95;
  output c0sm_b0m_v0m_n120;
  output c0sm_b0m_v0m_n121;

  // moduleNum: x82
  // type: nor2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1483/1488
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:252 c0sm_b0m_v0m_n120 c0sm_b0m_v0m_n121 
  // group: sel; nodes: [ c0sm_b0m_n2 ]

  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u187 (.A(c0sm_b0m_v0m_n94), .B(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n121));
  NOR2_X0P5A_A12TR c0sm_b0m_v0m_u185 (.A(c0sm_b0m_v0m_n95), .B(c0sm_b0m_n2), .Y(c0sm_b0m_v0m_n120));
endmodule
module nor2gate_mx83 
(
  c0sm_n3, 
  c0sm_v0m_n9, 
  reset, 
  c0sm_b0m_n9,
  c0sm_v0m_n13
);
  input c0sm_n3;
  input c0sm_v0m_n9;
  input reset;
  output c0sm_b0m_n9;
  output c0sm_v0m_n13;
  wire debitout_1;

  // moduleNum: x83
  // type: nor2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 3
  // number of non-inferred gates: 0
  // ILP vars: 1492/1496
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:253 c0sm_v0m_n13 c0sm_b0m_n9 
  // group: sel; nodes: [ c0sm_v0m_n9 ]

  NOR2B_X0P5M_A12TR c0sm_b0m_u27 (.AN(debitout_1), .B(reset), .Y(c0sm_b0m_n9));
  NOR2_X0P5A_A12TR c0sm_v0m_u30 (.A(c0sm_v0m_n9), .B(c0sm_n3), .Y(c0sm_v0m_n13));
  INV_X0P5B_A12TR c0sm_v0m_u10 (.A(c0sm_v0m_n9), .Y(debitout_1));
endmodule
module nor2gate_mx84 
(
  c0sm_v0m_n1, 
  c0sm_v0m_n2, 
  c0sm_v0m_n6, 
  c0sm_v0m_n32,
  c0sm_v0m_n33
);
  input c0sm_v0m_n1;
  input c0sm_v0m_n2;
  input c0sm_v0m_n6;
  output c0sm_v0m_n32;
  output c0sm_v0m_n33;

  // moduleNum: x84
  // type: nor2gate
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 0
  // number of word inputs: 0
  // number of word outputs: 1
  // number of internal gates: 2
  // number of non-inferred gates: 0
  // ILP vars: 1501/1501
  // type: INFERRED
  // marked bad? no
  // output word of size 2 : index:236 c0sm_v0m_n32 c0sm_v0m_n33 
  // group: sel; nodes: [ c0sm_v0m_n1 ]

  NOR2_X0P5A_A12TR c0sm_v0m_u6 (.A(c0sm_v0m_n1), .B(c0sm_v0m_n6), .Y(c0sm_v0m_n33));
  NOR2_X0P5A_A12TR c0sm_v0m_u3 (.A(c0sm_v0m_n1), .B(c0sm_v0m_n2), .Y(c0sm_v0m_n32));
endmodule
module mux_merged_mx85 
(
  c0nm_b0m_v0m_n105, 
  c0nm_b0m_v0m_n107, 
  c0nm_b0m_v0m_n108, 
  c0nm_b0m_v0m_n109, 
  c0nm_b0m_v0m_n122, 
  c0nm_b0m_v0m_n25, 
  c0nm_b0m_v0m_n27, 
  c0nm_b0m_v0m_n31, 
  c0nm_b0m_v0m_n32, 
  reset, 
  c0nm_b0m_v0m_n218,
  c0nm_b0m_v0m_n219
);
  input c0nm_b0m_v0m_n105;
  input c0nm_b0m_v0m_n107;
  input c0nm_b0m_v0m_n108;
  input c0nm_b0m_v0m_n109;
  input c0nm_b0m_v0m_n122;
  input c0nm_b0m_v0m_n25;
  input c0nm_b0m_v0m_n27;
  input c0nm_b0m_v0m_n31;
  input c0nm_b0m_v0m_n32;
  input reset;
  output c0nm_b0m_v0m_n218;
  output c0nm_b0m_v0m_n219;
  wire c0nm_b0m_v0m_n106;
  wire c0nm_b0m_v0m_n123;

  // moduleNum: x85
  // type: mux_merged
  // conflicting modules: 
  // number of bit inputs: 10
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 4
  // number of non-inferred gates: 0
  // ILP vars: 1518/1520
  // type: INFERRED
  // marked bad? no
  // merged: mux21i_mx11 mux21i_aoi221_mx112 mux21i_aoi221_mx114 mux21i_aoi221_mx157 
  // group: sel; nodes: [ c0nm_b0m_v0m_n107 reset c0nm_b0m_v0m_n108 c0nm_b0m_v0m_n109 ]

  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u92 (.A0(c0nm_b0m_v0m_n108), .A1(c0nm_b0m_v0m_n31), .B0(c0nm_b0m_v0m_n109), .B1(c0nm_b0m_v0m_n32), .C0(reset), .Y(c0nm_b0m_v0m_n123));
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u91 (.A(c0nm_b0m_v0m_n122), .B(c0nm_b0m_v0m_n123), .S0(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n218));
  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u85 (.A0(c0nm_b0m_v0m_n108), .A1(c0nm_b0m_v0m_n25), .B0(c0nm_b0m_v0m_n109), .B1(c0nm_b0m_v0m_n27), .C0(reset), .Y(c0nm_b0m_v0m_n106));
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u84 (.A(c0nm_b0m_v0m_n105), .B(c0nm_b0m_v0m_n106), .S0(c0nm_b0m_v0m_n107), .Y(c0nm_b0m_v0m_n219));
endmodule
module mux_merged_mx86 
(
  c0nm_b0m_v0m_n25, 
  c0nm_b0m_v0m_n27, 
  c0nm_b0m_v0m_n31, 
  c0nm_b0m_v0m_n32, 
  c0nm_b0m_v0m_n74, 
  c0nm_b0m_v0m_n76, 
  c0nm_b0m_v0m_n77, 
  c0nm_b0m_v0m_n78, 
  c0nm_b0m_v0m_n79, 
  reset, 
  c0nm_b0m_v0m_n242,
  c0nm_b0m_v0m_n243
);
  input c0nm_b0m_v0m_n25;
  input c0nm_b0m_v0m_n27;
  input c0nm_b0m_v0m_n31;
  input c0nm_b0m_v0m_n32;
  input c0nm_b0m_v0m_n74;
  input c0nm_b0m_v0m_n76;
  input c0nm_b0m_v0m_n77;
  input c0nm_b0m_v0m_n78;
  input c0nm_b0m_v0m_n79;
  input reset;
  output c0nm_b0m_v0m_n242;
  output c0nm_b0m_v0m_n243;
  wire c0nm_b0m_v0m_n75;
  wire c0nm_b0m_v0m_n80;

  // moduleNum: x86
  // type: mux_merged
  // conflicting modules: 
  // number of bit inputs: 10
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 4
  // number of non-inferred gates: 0
  // ILP vars: 1524/1526
  // type: INFERRED
  // marked bad? no
  // merged: mux21i_mx13 mux21i_aoi221_mx121 mux21i_aoi221_mx122 mux21i_aoi221_mx168 
  // group: sel; nodes: [ c0nm_b0m_v0m_n76 reset c0nm_b0m_v0m_n77 c0nm_b0m_v0m_n78 ]

  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u38 (.A0(c0nm_b0m_v0m_n77), .A1(c0nm_b0m_v0m_n31), .B0(c0nm_b0m_v0m_n78), .B1(c0nm_b0m_v0m_n32), .C0(reset), .Y(c0nm_b0m_v0m_n80));
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u37 (.A(c0nm_b0m_v0m_n79), .B(c0nm_b0m_v0m_n80), .S0(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n242));
  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u35 (.A0(c0nm_b0m_v0m_n77), .A1(c0nm_b0m_v0m_n25), .B0(c0nm_b0m_v0m_n78), .B1(c0nm_b0m_v0m_n27), .C0(reset), .Y(c0nm_b0m_v0m_n75));
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u34 (.A(c0nm_b0m_v0m_n74), .B(c0nm_b0m_v0m_n75), .S0(c0nm_b0m_v0m_n76), .Y(c0nm_b0m_v0m_n243));
endmodule
module mux_merged_mx87 
(
  c0nm_b0m_v0m_n22, 
  c0nm_b0m_v0m_n23, 
  c0nm_b0m_v0m_n25, 
  c0nm_b0m_v0m_n26, 
  c0nm_b0m_v0m_n27, 
  c0nm_b0m_v0m_n28, 
  c0nm_b0m_v0m_n29, 
  c0nm_b0m_v0m_n31, 
  c0nm_b0m_v0m_n32, 
  reset, 
  c0nm_b0m_v0m_n253,
  c0nm_b0m_v0m_n254
);
  input c0nm_b0m_v0m_n22;
  input c0nm_b0m_v0m_n23;
  input c0nm_b0m_v0m_n25;
  input c0nm_b0m_v0m_n26;
  input c0nm_b0m_v0m_n27;
  input c0nm_b0m_v0m_n28;
  input c0nm_b0m_v0m_n29;
  input c0nm_b0m_v0m_n31;
  input c0nm_b0m_v0m_n32;
  input reset;
  output c0nm_b0m_v0m_n253;
  output c0nm_b0m_v0m_n254;
  wire c0nm_b0m_v0m_n24;
  wire c0nm_b0m_v0m_n30;

  // moduleNum: x87
  // type: mux_merged
  // conflicting modules: 
  // number of bit inputs: 10
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 4
  // number of non-inferred gates: 0
  // ILP vars: 1527/1529
  // type: INFERRED
  // marked bad? no
  // merged: mux21i_mx14 mux21i_aoi221_mx111 mux21i_aoi221_mx113 mux21i_aoi221_mx156 
  // group: sel; nodes: [ c0nm_b0m_v0m_n22 reset c0nm_b0m_v0m_n28 c0nm_b0m_v0m_n26 ]

  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u21 (.A0(c0nm_b0m_v0m_n31), .A1(c0nm_b0m_v0m_n26), .B0(c0nm_b0m_v0m_n32), .B1(c0nm_b0m_v0m_n28), .C0(reset), .Y(c0nm_b0m_v0m_n30));
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u20 (.A(c0nm_b0m_v0m_n29), .B(c0nm_b0m_v0m_n30), .S0(c0nm_b0m_v0m_n22), .Y(c0nm_b0m_v0m_n253));
  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u19 (.A0(c0nm_b0m_v0m_n25), .A1(c0nm_b0m_v0m_n26), .B0(c0nm_b0m_v0m_n27), .B1(c0nm_b0m_v0m_n28), .C0(reset), .Y(c0nm_b0m_v0m_n24));
  MXIT2_X0P5M_A12TR c0nm_b0m_v0m_u18 (.A(c0nm_b0m_v0m_n23), .B(c0nm_b0m_v0m_n24), .S0(c0nm_b0m_v0m_n22), .Y(c0nm_b0m_v0m_n254));
endmodule
module mux_merged_mx88 
(
  c0sm_b0m_v0m_n105, 
  c0sm_b0m_v0m_n107, 
  c0sm_b0m_v0m_n108, 
  c0sm_b0m_v0m_n109, 
  c0sm_b0m_v0m_n122, 
  c0sm_b0m_v0m_n25, 
  c0sm_b0m_v0m_n27, 
  c0sm_b0m_v0m_n31, 
  c0sm_b0m_v0m_n32, 
  reset, 
  c0sm_b0m_v0m_n319,
  c0sm_b0m_v0m_n320
);
  input c0sm_b0m_v0m_n105;
  input c0sm_b0m_v0m_n107;
  input c0sm_b0m_v0m_n108;
  input c0sm_b0m_v0m_n109;
  input c0sm_b0m_v0m_n122;
  input c0sm_b0m_v0m_n25;
  input c0sm_b0m_v0m_n27;
  input c0sm_b0m_v0m_n31;
  input c0sm_b0m_v0m_n32;
  input reset;
  output c0sm_b0m_v0m_n319;
  output c0sm_b0m_v0m_n320;
  wire c0sm_b0m_v0m_n106;
  wire c0sm_b0m_v0m_n123;

  // moduleNum: x88
  // type: mux_merged
  // conflicting modules: 
  // number of bit inputs: 10
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 4
  // number of non-inferred gates: 0
  // ILP vars: 1530/1532
  // type: INFERRED
  // marked bad? no
  // merged: mux21i_mx17 mux21i_aoi221_mx124 mux21i_aoi221_mx126 mux21i_aoi221_mx193 
  // group: sel; nodes: [ c0sm_b0m_v0m_n107 reset c0sm_b0m_v0m_n108 c0sm_b0m_v0m_n109 ]

  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u92 (.A0(c0sm_b0m_v0m_n108), .A1(c0sm_b0m_v0m_n31), .B0(c0sm_b0m_v0m_n109), .B1(c0sm_b0m_v0m_n32), .C0(reset), .Y(c0sm_b0m_v0m_n123));
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u91 (.A(c0sm_b0m_v0m_n122), .B(c0sm_b0m_v0m_n123), .S0(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n320));
  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u85 (.A0(c0sm_b0m_v0m_n108), .A1(c0sm_b0m_v0m_n25), .B0(c0sm_b0m_v0m_n109), .B1(c0sm_b0m_v0m_n27), .C0(reset), .Y(c0sm_b0m_v0m_n106));
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u84 (.A(c0sm_b0m_v0m_n105), .B(c0sm_b0m_v0m_n106), .S0(c0sm_b0m_v0m_n107), .Y(c0sm_b0m_v0m_n319));
endmodule
module mux_merged_mx89 
(
  c0sm_b0m_v0m_n25, 
  c0sm_b0m_v0m_n27, 
  c0sm_b0m_v0m_n31, 
  c0sm_b0m_v0m_n32, 
  c0sm_b0m_v0m_n74, 
  c0sm_b0m_v0m_n76, 
  c0sm_b0m_v0m_n77, 
  c0sm_b0m_v0m_n78, 
  c0sm_b0m_v0m_n79, 
  reset, 
  c0sm_b0m_v0m_n295,
  c0sm_b0m_v0m_n296
);
  input c0sm_b0m_v0m_n25;
  input c0sm_b0m_v0m_n27;
  input c0sm_b0m_v0m_n31;
  input c0sm_b0m_v0m_n32;
  input c0sm_b0m_v0m_n74;
  input c0sm_b0m_v0m_n76;
  input c0sm_b0m_v0m_n77;
  input c0sm_b0m_v0m_n78;
  input c0sm_b0m_v0m_n79;
  input reset;
  output c0sm_b0m_v0m_n295;
  output c0sm_b0m_v0m_n296;
  wire c0sm_b0m_v0m_n75;
  wire c0sm_b0m_v0m_n80;

  // moduleNum: x89
  // type: mux_merged
  // conflicting modules: 
  // number of bit inputs: 10
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 4
  // number of non-inferred gates: 0
  // ILP vars: 1536/1538
  // type: INFERRED
  // marked bad? no
  // merged: mux21i_mx19 mux21i_aoi221_mx133 mux21i_aoi221_mx134 mux21i_aoi221_mx204 
  // group: sel; nodes: [ c0sm_b0m_v0m_n76 reset c0sm_b0m_v0m_n77 c0sm_b0m_v0m_n78 ]

  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u38 (.A0(c0sm_b0m_v0m_n77), .A1(c0sm_b0m_v0m_n31), .B0(c0sm_b0m_v0m_n78), .B1(c0sm_b0m_v0m_n32), .C0(reset), .Y(c0sm_b0m_v0m_n80));
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u37 (.A(c0sm_b0m_v0m_n79), .B(c0sm_b0m_v0m_n80), .S0(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n296));
  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u35 (.A0(c0sm_b0m_v0m_n77), .A1(c0sm_b0m_v0m_n25), .B0(c0sm_b0m_v0m_n78), .B1(c0sm_b0m_v0m_n27), .C0(reset), .Y(c0sm_b0m_v0m_n75));
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u34 (.A(c0sm_b0m_v0m_n74), .B(c0sm_b0m_v0m_n75), .S0(c0sm_b0m_v0m_n76), .Y(c0sm_b0m_v0m_n295));
endmodule
module mux_merged_mx90 
(
  c0sm_b0m_v0m_n22, 
  c0sm_b0m_v0m_n23, 
  c0sm_b0m_v0m_n25, 
  c0sm_b0m_v0m_n26, 
  c0sm_b0m_v0m_n27, 
  c0sm_b0m_v0m_n28, 
  c0sm_b0m_v0m_n29, 
  c0sm_b0m_v0m_n31, 
  c0sm_b0m_v0m_n32, 
  reset, 
  c0sm_b0m_v0m_n284,
  c0sm_b0m_v0m_n285
);
  input c0sm_b0m_v0m_n22;
  input c0sm_b0m_v0m_n23;
  input c0sm_b0m_v0m_n25;
  input c0sm_b0m_v0m_n26;
  input c0sm_b0m_v0m_n27;
  input c0sm_b0m_v0m_n28;
  input c0sm_b0m_v0m_n29;
  input c0sm_b0m_v0m_n31;
  input c0sm_b0m_v0m_n32;
  input reset;
  output c0sm_b0m_v0m_n284;
  output c0sm_b0m_v0m_n285;
  wire c0sm_b0m_v0m_n24;
  wire c0sm_b0m_v0m_n30;

  // moduleNum: x90
  // type: mux_merged
  // conflicting modules: 
  // number of bit inputs: 10
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 4
  // number of non-inferred gates: 0
  // ILP vars: 1539/1541
  // type: INFERRED
  // marked bad? no
  // merged: mux21i_mx20 mux21i_aoi221_mx123 mux21i_aoi221_mx125 mux21i_aoi221_mx192 
  // group: sel; nodes: [ c0sm_b0m_v0m_n22 reset c0sm_b0m_v0m_n28 c0sm_b0m_v0m_n26 ]

  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u21 (.A0(c0sm_b0m_v0m_n31), .A1(c0sm_b0m_v0m_n26), .B0(c0sm_b0m_v0m_n32), .B1(c0sm_b0m_v0m_n28), .C0(reset), .Y(c0sm_b0m_v0m_n30));
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u20 (.A(c0sm_b0m_v0m_n29), .B(c0sm_b0m_v0m_n30), .S0(c0sm_b0m_v0m_n22), .Y(c0sm_b0m_v0m_n285));
  AOI221_X0P5M_A12TR c0sm_b0m_v0m_u19 (.A0(c0sm_b0m_v0m_n25), .A1(c0sm_b0m_v0m_n26), .B0(c0sm_b0m_v0m_n27), .B1(c0sm_b0m_v0m_n28), .C0(reset), .Y(c0sm_b0m_v0m_n24));
  MXIT2_X0P5M_A12TR c0sm_b0m_v0m_u18 (.A(c0sm_b0m_v0m_n23), .B(c0sm_b0m_v0m_n24), .S0(c0sm_b0m_v0m_n22), .Y(c0sm_b0m_v0m_n284));
endmodule
module mux_merged_mx91 
(
  c0nm_b0m_v0m_buffers0_10_, 
  c0nm_b0m_v0m_buffers0_11_, 
  c0nm_b0m_v0m_buffers0_2_, 
  c0nm_b0m_v0m_buffers0_4_, 
  c0nm_b0m_v0m_buffers0_7_, 
  c0nm_b0m_v0m_buffers0_8_, 
  c0nm_b0m_v0m_buffers0_9_, 
  c0nm_b0m_v0m_n131, 
  c0nm_b0m_v0m_n134, 
  c0nm_b0m_v0m_n144, 
  c0nm_b0m_v0m_n147, 
  c0nm_b0m_v0m_n162, 
  c0nm_b0m_v0m_n165, 
  c0nm_b0m_v0m_n168, 
  c0nm_b0m_v0m_n171, 
  c0nm_b0m_v0m_n174, 
  c0nm_b0m_v0m_n177, 
  c0nm_b0m_v0m_n180, 
  c0nm_b0m_v0m_n183, 
  c0nm_b0m_v0m_n186, 
  c0nm_b0m_v0m_n187, 
  c0nm_b0m_v0m_n190, 
  c0nm_b0m_v0m_n192, 
  c0nm_b0m_v0m_n193, 
  c0nm_b0m_v0m_n21, 
  c0nm_b0m_v0m_n35, 
  c0nm_b0m_v0m_n41, 
  c0nm_b0m_v0m_n62, 
  c0nm_b0m_v0m_n65, 
  c0nm_b0m_v0m_n68, 
  c0nm_b0m_v0m_n71, 
  c0nm_b0m_v0m_n73, 
  c0nm_b0m_headflit_10_,
  c0nm_b0m_headflit_11_,
  c0nm_b0m_headflit_8_,
  c0nm_b0m_headflit_9_,
  c0nm_headflit_2_,
  c0nm_headflit_4_,
  c0nm_headflit_7_
);
  input c0nm_b0m_v0m_buffers0_10_;
  input c0nm_b0m_v0m_buffers0_11_;
  input c0nm_b0m_v0m_buffers0_2_;
  input c0nm_b0m_v0m_buffers0_4_;
  input c0nm_b0m_v0m_buffers0_7_;
  input c0nm_b0m_v0m_buffers0_8_;
  input c0nm_b0m_v0m_buffers0_9_;
  input c0nm_b0m_v0m_n131;
  input c0nm_b0m_v0m_n134;
  input c0nm_b0m_v0m_n144;
  input c0nm_b0m_v0m_n147;
  input c0nm_b0m_v0m_n162;
  input c0nm_b0m_v0m_n165;
  input c0nm_b0m_v0m_n168;
  input c0nm_b0m_v0m_n171;
  input c0nm_b0m_v0m_n174;
  input c0nm_b0m_v0m_n177;
  input c0nm_b0m_v0m_n180;
  input c0nm_b0m_v0m_n183;
  input c0nm_b0m_v0m_n186;
  input c0nm_b0m_v0m_n187;
  input c0nm_b0m_v0m_n190;
  input c0nm_b0m_v0m_n192;
  input c0nm_b0m_v0m_n193;
  input c0nm_b0m_v0m_n21;
  input c0nm_b0m_v0m_n35;
  input c0nm_b0m_v0m_n41;
  input c0nm_b0m_v0m_n62;
  input c0nm_b0m_v0m_n65;
  input c0nm_b0m_v0m_n68;
  input c0nm_b0m_v0m_n71;
  input c0nm_b0m_v0m_n73;
  output c0nm_b0m_headflit_10_;
  output c0nm_b0m_headflit_11_;
  output c0nm_b0m_headflit_8_;
  output c0nm_b0m_headflit_9_;
  output c0nm_headflit_2_;
  output c0nm_headflit_4_;
  output c0nm_headflit_7_;
  wire c0nm_b0m_v0m_n265;
  wire c0nm_b0m_v0m_n266;
  wire c0nm_b0m_v0m_n267;
  wire c0nm_b0m_v0m_n270;
  wire c0nm_b0m_v0m_n272;
  wire c0nm_b0m_v0m_n273;
  wire c0nm_b0m_v0m_n274;

  // moduleNum: x91
  // type: mux_merged
  // conflicting modules: 
  // number of bit inputs: 32
  // number of bit outputs: 7
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 14
  // number of non-inferred gates: 0
  // ILP vars: 1542/1554
  // type: INFERRED
  // marked bad? no
  // merged: mux21i_aoi22_mx42 mux21i_oai221_mx217 
  // group: sel; nodes: [ c0nm_b0m_v0m_n193 c0nm_b0m_v0m_n192 c0nm_b0m_v0m_n187 c0nm_b0m_v0m_n73 ]

  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u256 (.A0(c0nm_b0m_v0m_buffers0_10_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n183), .Y(c0nm_b0m_v0m_n274));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u255 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n180), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n71), .C0(c0nm_b0m_v0m_n274), .Y(c0nm_b0m_headflit_10_));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u251 (.A0(c0nm_b0m_v0m_n193), .A1(c0nm_b0m_v0m_buffers0_11_), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n190), .Y(c0nm_b0m_v0m_n273));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u250 (.A0(c0nm_b0m_v0m_n186), .A1(c0nm_b0m_v0m_n187), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n21), .C0(c0nm_b0m_v0m_n273), .Y(c0nm_b0m_headflit_11_));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u246 (.A0(c0nm_b0m_v0m_buffers0_2_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n134), .Y(c0nm_b0m_v0m_n272));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u245 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n131), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n35), .C0(c0nm_b0m_v0m_n272), .Y(c0nm_headflit_2_));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u236 (.A0(c0nm_b0m_v0m_buffers0_4_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n147), .Y(c0nm_b0m_v0m_n270));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u235 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n144), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n41), .C0(c0nm_b0m_v0m_n270), .Y(c0nm_headflit_4_));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u221 (.A0(c0nm_b0m_v0m_buffers0_7_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n165), .Y(c0nm_b0m_v0m_n267));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u220 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n162), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n62), .C0(c0nm_b0m_v0m_n267), .Y(c0nm_headflit_7_));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u216 (.A0(c0nm_b0m_v0m_buffers0_8_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n171), .Y(c0nm_b0m_v0m_n266));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u215 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n168), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n65), .C0(c0nm_b0m_v0m_n266), .Y(c0nm_b0m_headflit_8_));
  AOI22_X0P5M_A12TR c0nm_b0m_v0m_u211 (.A0(c0nm_b0m_v0m_buffers0_9_), .A1(c0nm_b0m_v0m_n193), .B0(c0nm_b0m_v0m_n192), .B1(c0nm_b0m_v0m_n177), .Y(c0nm_b0m_v0m_n265));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u210 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n174), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n68), .C0(c0nm_b0m_v0m_n265), .Y(c0nm_b0m_headflit_9_));
endmodule
module mux_merged_mx92 
(
  c0sm_b0m_v0m_buffers0_0_, 
  c0sm_b0m_v0m_buffers0_10_, 
  c0sm_b0m_v0m_buffers0_11_, 
  c0sm_b0m_v0m_buffers0_1_, 
  c0sm_b0m_v0m_buffers0_2_, 
  c0sm_b0m_v0m_buffers0_4_, 
  c0sm_b0m_v0m_buffers0_7_, 
  c0sm_b0m_v0m_buffers0_8_, 
  c0sm_b0m_v0m_buffers0_9_, 
  c0sm_b0m_v0m_n105, 
  c0sm_b0m_v0m_n114, 
  c0sm_b0m_v0m_n122, 
  c0sm_b0m_v0m_n125, 
  c0sm_b0m_v0m_n131, 
  c0sm_b0m_v0m_n134, 
  c0sm_b0m_v0m_n144, 
  c0sm_b0m_v0m_n147, 
  c0sm_b0m_v0m_n162, 
  c0sm_b0m_v0m_n165, 
  c0sm_b0m_v0m_n168, 
  c0sm_b0m_v0m_n171, 
  c0sm_b0m_v0m_n174, 
  c0sm_b0m_v0m_n177, 
  c0sm_b0m_v0m_n180, 
  c0sm_b0m_v0m_n183, 
  c0sm_b0m_v0m_n186, 
  c0sm_b0m_v0m_n187, 
  c0sm_b0m_v0m_n190, 
  c0sm_b0m_v0m_n192, 
  c0sm_b0m_v0m_n193, 
  c0sm_b0m_v0m_n21, 
  c0sm_b0m_v0m_n23, 
  c0sm_b0m_v0m_n29, 
  c0sm_b0m_v0m_n35, 
  c0sm_b0m_v0m_n41, 
  c0sm_b0m_v0m_n62, 
  c0sm_b0m_v0m_n65, 
  c0sm_b0m_v0m_n68, 
  c0sm_b0m_v0m_n71, 
  c0sm_b0m_v0m_n73, 
  c0sm_b0m_headflit_10_,
  c0sm_b0m_headflit_11_,
  c0sm_b0m_headflit_8_,
  c0sm_b0m_headflit_9_,
  c0sm_headflit_0_,
  c0sm_headflit_1_,
  c0sm_headflit_2_,
  c0sm_headflit_4_,
  c0sm_headflit_7_
);
  input c0sm_b0m_v0m_buffers0_0_;
  input c0sm_b0m_v0m_buffers0_10_;
  input c0sm_b0m_v0m_buffers0_11_;
  input c0sm_b0m_v0m_buffers0_1_;
  input c0sm_b0m_v0m_buffers0_2_;
  input c0sm_b0m_v0m_buffers0_4_;
  input c0sm_b0m_v0m_buffers0_7_;
  input c0sm_b0m_v0m_buffers0_8_;
  input c0sm_b0m_v0m_buffers0_9_;
  input c0sm_b0m_v0m_n105;
  input c0sm_b0m_v0m_n114;
  input c0sm_b0m_v0m_n122;
  input c0sm_b0m_v0m_n125;
  input c0sm_b0m_v0m_n131;
  input c0sm_b0m_v0m_n134;
  input c0sm_b0m_v0m_n144;
  input c0sm_b0m_v0m_n147;
  input c0sm_b0m_v0m_n162;
  input c0sm_b0m_v0m_n165;
  input c0sm_b0m_v0m_n168;
  input c0sm_b0m_v0m_n171;
  input c0sm_b0m_v0m_n174;
  input c0sm_b0m_v0m_n177;
  input c0sm_b0m_v0m_n180;
  input c0sm_b0m_v0m_n183;
  input c0sm_b0m_v0m_n186;
  input c0sm_b0m_v0m_n187;
  input c0sm_b0m_v0m_n190;
  input c0sm_b0m_v0m_n192;
  input c0sm_b0m_v0m_n193;
  input c0sm_b0m_v0m_n21;
  input c0sm_b0m_v0m_n23;
  input c0sm_b0m_v0m_n29;
  input c0sm_b0m_v0m_n35;
  input c0sm_b0m_v0m_n41;
  input c0sm_b0m_v0m_n62;
  input c0sm_b0m_v0m_n65;
  input c0sm_b0m_v0m_n68;
  input c0sm_b0m_v0m_n71;
  input c0sm_b0m_v0m_n73;
  output c0sm_b0m_headflit_10_;
  output c0sm_b0m_headflit_11_;
  output c0sm_b0m_headflit_8_;
  output c0sm_b0m_headflit_9_;
  output c0sm_headflit_0_;
  output c0sm_headflit_1_;
  output c0sm_headflit_2_;
  output c0sm_headflit_4_;
  output c0sm_headflit_7_;
  wire c0sm_b0m_v0m_n265;
  wire c0sm_b0m_v0m_n266;
  wire c0sm_b0m_v0m_n267;
  wire c0sm_b0m_v0m_n270;
  wire c0sm_b0m_v0m_n272;
  wire c0sm_b0m_v0m_n273;
  wire c0sm_b0m_v0m_n274;
  wire c0sm_b0m_v0m_n275;
  wire c0sm_b0m_v0m_n276;

  // moduleNum: x92
  // type: mux_merged
  // conflicting modules: 
  // number of bit inputs: 40
  // number of bit outputs: 9
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 18
  // number of non-inferred gates: 0
  // ILP vars: 1605/1617
  // type: INFERRED
  // marked bad? no
  // merged: mux21i_aoi22_mx77 mux21i_oai221_mx231 
  // group: sel; nodes: [ c0sm_b0m_v0m_n193 c0sm_b0m_v0m_n192 c0sm_b0m_v0m_n187 c0sm_b0m_v0m_n73 ]

  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u269 (.A0(c0sm_b0m_v0m_buffers0_0_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n114), .Y(c0sm_b0m_v0m_n276));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u268 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n105), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n23), .C0(c0sm_b0m_v0m_n276), .Y(c0sm_headflit_0_));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u264 (.A0(c0sm_b0m_v0m_buffers0_1_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n125), .Y(c0sm_b0m_v0m_n275));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u263 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n122), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n29), .C0(c0sm_b0m_v0m_n275), .Y(c0sm_headflit_1_));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u256 (.A0(c0sm_b0m_v0m_buffers0_10_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n183), .Y(c0sm_b0m_v0m_n274));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u255 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n180), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n71), .C0(c0sm_b0m_v0m_n274), .Y(c0sm_b0m_headflit_10_));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u251 (.A0(c0sm_b0m_v0m_n193), .A1(c0sm_b0m_v0m_buffers0_11_), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n190), .Y(c0sm_b0m_v0m_n273));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u250 (.A0(c0sm_b0m_v0m_n186), .A1(c0sm_b0m_v0m_n187), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n21), .C0(c0sm_b0m_v0m_n273), .Y(c0sm_b0m_headflit_11_));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u246 (.A0(c0sm_b0m_v0m_buffers0_2_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n134), .Y(c0sm_b0m_v0m_n272));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u245 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n131), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n35), .C0(c0sm_b0m_v0m_n272), .Y(c0sm_headflit_2_));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u236 (.A0(c0sm_b0m_v0m_buffers0_4_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n147), .Y(c0sm_b0m_v0m_n270));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u235 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n144), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n41), .C0(c0sm_b0m_v0m_n270), .Y(c0sm_headflit_4_));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u221 (.A0(c0sm_b0m_v0m_buffers0_7_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n165), .Y(c0sm_b0m_v0m_n267));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u220 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n162), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n62), .C0(c0sm_b0m_v0m_n267), .Y(c0sm_headflit_7_));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u216 (.A0(c0sm_b0m_v0m_buffers0_8_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n171), .Y(c0sm_b0m_v0m_n266));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u215 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n168), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n65), .C0(c0sm_b0m_v0m_n266), .Y(c0sm_b0m_headflit_8_));
  AOI22_X0P5M_A12TR c0sm_b0m_v0m_u211 (.A0(c0sm_b0m_v0m_buffers0_9_), .A1(c0sm_b0m_v0m_n193), .B0(c0sm_b0m_v0m_n192), .B1(c0sm_b0m_v0m_n177), .Y(c0sm_b0m_v0m_n265));
  OAI221_X0P5M_A12TR c0sm_b0m_v0m_u210 (.A0(c0sm_b0m_v0m_n187), .A1(c0sm_b0m_v0m_n174), .B0(c0sm_b0m_v0m_n73), .B1(c0sm_b0m_v0m_n68), .C0(c0sm_b0m_v0m_n265), .Y(c0sm_b0m_headflit_9_));
endmodule
module mux_merged_mx93 
(
  c0nm_b0m_v0m_buffers0_0_, 
  c0nm_b0m_v0m_n105, 
  c0nm_b0m_v0m_n110, 
  c0nm_b0m_v0m_n111, 
  c0nm_b0m_v0m_n113, 
  c0nm_b0m_v0m_n114, 
  c0nm_b0m_v0m_n115, 
  c0nm_b0m_v0m_n187, 
  c0nm_b0m_v0m_n192, 
  c0nm_b0m_v0m_n193, 
  c0nm_b0m_v0m_n23, 
  c0nm_b0m_v0m_n276, 
  c0nm_b0m_v0m_n73, 
  debitout_0, 
  c0nm_b0m_v0m_n27,
  c0nm_headflit_0_
);
  input c0nm_b0m_v0m_buffers0_0_;
  input c0nm_b0m_v0m_n105;
  input c0nm_b0m_v0m_n110;
  input c0nm_b0m_v0m_n111;
  input c0nm_b0m_v0m_n113;
  input c0nm_b0m_v0m_n114;
  input c0nm_b0m_v0m_n115;
  input c0nm_b0m_v0m_n187;
  input c0nm_b0m_v0m_n192;
  input c0nm_b0m_v0m_n193;
  input c0nm_b0m_v0m_n23;
  input c0nm_b0m_v0m_n276;
  input c0nm_b0m_v0m_n73;
  input debitout_0;
  output c0nm_b0m_v0m_n27;
  output c0nm_headflit_0_;
  wire c0nm_b0m_v0m_n112;

  // moduleNum: x93
  // type: mux_merged
  // conflicting modules: 
  // number of bit inputs: 14
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 3
  // number of non-inferred gates: 0
  // ILP vars: 1668/1668
  // type: INFERRED
  // marked bad? no
  // merged: mux21i_aoi221_mx136 mux21i_aoi221_mx139 mux21i_aoi221_mx142 mux21i_aoi221_mx145 mux21i_aoi221_mx148
  // mux21i_aoi221_mx149 mux21i_aoi221_mx159 mux21i_aoi221_mx162 mux21i_oai221_mx218
  // group: sel; nodes: [ c0nm_b0m_v0m_n193 c0nm_b0m_v0m_n114 c0nm_b0m_v0m_buffers0_0_ c0nm_b0m_v0m_n192 c0nm_b0m_v0m_n115
  // c0nm_b0m_v0m_n113 c0nm_b0m_v0m_n105 c0nm_b0m_v0m_n23 ]

  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u268 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n105), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n23), .C0(c0nm_b0m_v0m_n276), .Y(c0nm_headflit_0_));
  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u87 (.A0(c0nm_b0m_v0m_n113), .A1(c0nm_b0m_v0m_n114), .B0(c0nm_b0m_v0m_buffers0_0_), .B1(c0nm_b0m_v0m_n115), .C0(debitout_0), .Y(c0nm_b0m_v0m_n112));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u86 (.A0(c0nm_b0m_v0m_n110), .A1(c0nm_b0m_v0m_n105), .B0(c0nm_b0m_v0m_n111), .B1(c0nm_b0m_v0m_n23), .C0(c0nm_b0m_v0m_n112), .Y(c0nm_b0m_v0m_n27));
endmodule
module mux_merged_mx94 
(
  c0nm_b0m_v0m_buffers0_1_, 
  c0nm_b0m_v0m_n110, 
  c0nm_b0m_v0m_n111, 
  c0nm_b0m_v0m_n113, 
  c0nm_b0m_v0m_n115, 
  c0nm_b0m_v0m_n122, 
  c0nm_b0m_v0m_n125, 
  c0nm_b0m_v0m_n187, 
  c0nm_b0m_v0m_n192, 
  c0nm_b0m_v0m_n193, 
  c0nm_b0m_v0m_n275, 
  c0nm_b0m_v0m_n29, 
  c0nm_b0m_v0m_n73, 
  debitout_0, 
  c0nm_b0m_v0m_n32,
  c0nm_headflit_1_
);
  input c0nm_b0m_v0m_buffers0_1_;
  input c0nm_b0m_v0m_n110;
  input c0nm_b0m_v0m_n111;
  input c0nm_b0m_v0m_n113;
  input c0nm_b0m_v0m_n115;
  input c0nm_b0m_v0m_n122;
  input c0nm_b0m_v0m_n125;
  input c0nm_b0m_v0m_n187;
  input c0nm_b0m_v0m_n192;
  input c0nm_b0m_v0m_n193;
  input c0nm_b0m_v0m_n275;
  input c0nm_b0m_v0m_n29;
  input c0nm_b0m_v0m_n73;
  input debitout_0;
  output c0nm_b0m_v0m_n32;
  output c0nm_headflit_1_;
  wire c0nm_b0m_v0m_n124;

  // moduleNum: x94
  // type: mux_merged
  // conflicting modules: 
  // number of bit inputs: 14
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 3
  // number of non-inferred gates: 0
  // ILP vars: 1669/1669
  // type: INFERRED
  // marked bad? no
  // merged: mux21i_aoi221_mx137 mux21i_aoi221_mx140 mux21i_aoi221_mx143 mux21i_aoi221_mx146 mux21i_aoi221_mx152
  // mux21i_aoi221_mx153 mux21i_aoi221_mx160 mux21i_aoi221_mx163 mux21i_oai221_mx219
  // group: sel; nodes: [ c0nm_b0m_v0m_n193 c0nm_b0m_v0m_n125 c0nm_b0m_v0m_buffers0_1_ c0nm_b0m_v0m_n192 c0nm_b0m_v0m_n115
  // c0nm_b0m_v0m_n113 c0nm_b0m_v0m_n122 c0nm_b0m_v0m_n29 ]

  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u263 (.A0(c0nm_b0m_v0m_n187), .A1(c0nm_b0m_v0m_n122), .B0(c0nm_b0m_v0m_n73), .B1(c0nm_b0m_v0m_n29), .C0(c0nm_b0m_v0m_n275), .Y(c0nm_headflit_1_));
  AOI221_X0P5M_A12TR c0nm_b0m_v0m_u94 (.A0(c0nm_b0m_v0m_n113), .A1(c0nm_b0m_v0m_n125), .B0(c0nm_b0m_v0m_buffers0_1_), .B1(c0nm_b0m_v0m_n115), .C0(debitout_0), .Y(c0nm_b0m_v0m_n124));
  OAI221_X0P5M_A12TR c0nm_b0m_v0m_u93 (.A0(c0nm_b0m_v0m_n110), .A1(c0nm_b0m_v0m_n122), .B0(c0nm_b0m_v0m_n111), .B1(c0nm_b0m_v0m_n29), .C0(c0nm_b0m_v0m_n124), .Y(c0nm_b0m_v0m_n32));
endmodule
module counter_mx95 
(
  c0nm_b0m_v0m_n257, 
  c0nm_b0m_v0m_n258, 
  clk, 
  c0nm_b0m_v0m_head_0_,
  c0nm_b0m_v0m_head_1_
);
  input c0nm_b0m_v0m_n257;
  input c0nm_b0m_v0m_n258;
  input clk;
  output c0nm_b0m_v0m_head_0_;
  output c0nm_b0m_v0m_head_1_;

  // moduleNum: x95
  // type: counter
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 4
  // number of non-inferred gates: 0
  // ILP vars: 1672/1672
  // type: INFERRED
  // marked bad? no

  DFFQ_X1M_A12TR c0nm_b0m_v0m_head_reg_1_ (.CK(clk), .Q(c0nm_b0m_v0m_head_1_), .D(c0nm_b0m_v0m_n257));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_head_reg_0_ (.CK(clk), .Q(c0nm_b0m_v0m_head_0_), .D(c0nm_b0m_v0m_n258));
endmodule
module counter_mx96 
(
  c0nm_b0m_v0m_n260, 
  c0nm_b0m_v0m_n261, 
  clk, 
  c0nm_b0m_v0m_tail_0_,
  c0nm_b0m_v0m_tail_1_
);
  input c0nm_b0m_v0m_n260;
  input c0nm_b0m_v0m_n261;
  input clk;
  output c0nm_b0m_v0m_tail_0_;
  output c0nm_b0m_v0m_tail_1_;

  // moduleNum: x96
  // type: counter
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 4
  // number of non-inferred gates: 0
  // ILP vars: 1673/1673
  // type: INFERRED
  // marked bad? no

  DFFQ_X1M_A12TR c0nm_b0m_v0m_tail_reg_0_ (.CK(clk), .Q(c0nm_b0m_v0m_tail_0_), .D(c0nm_b0m_v0m_n261));
  DFFQ_X1M_A12TR c0nm_b0m_v0m_tail_reg_1_ (.CK(clk), .Q(c0nm_b0m_v0m_tail_1_), .D(c0nm_b0m_v0m_n260));
endmodule
module counter_mx97 
(
  c0sm_b0m_v0m_n280, 
  c0sm_b0m_v0m_n281, 
  clk, 
  c0sm_b0m_v0m_head_0_,
  c0sm_b0m_v0m_head_1_
);
  input c0sm_b0m_v0m_n280;
  input c0sm_b0m_v0m_n281;
  input clk;
  output c0sm_b0m_v0m_head_0_;
  output c0sm_b0m_v0m_head_1_;

  // moduleNum: x97
  // type: counter
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 4
  // number of non-inferred gates: 0
  // ILP vars: 1674/1674
  // type: INFERRED
  // marked bad? no

  DFFQ_X1M_A12TR c0sm_b0m_v0m_head_reg_1_ (.CK(clk), .Q(c0sm_b0m_v0m_head_1_), .D(c0sm_b0m_v0m_n281));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_head_reg_0_ (.CK(clk), .Q(c0sm_b0m_v0m_head_0_), .D(c0sm_b0m_v0m_n280));
endmodule
module counter_mx98 
(
  c0sm_b0m_v0m_n277, 
  c0sm_b0m_v0m_n278, 
  clk, 
  c0sm_b0m_v0m_tail_0_,
  c0sm_b0m_v0m_tail_1_
);
  input c0sm_b0m_v0m_n277;
  input c0sm_b0m_v0m_n278;
  input clk;
  output c0sm_b0m_v0m_tail_0_;
  output c0sm_b0m_v0m_tail_1_;

  // moduleNum: x98
  // type: counter
  // conflicting modules: 
  // number of bit inputs: 3
  // number of bit outputs: 2
  // number of word inputs: 0
  // number of word outputs: 0
  // number of internal gates: 4
  // number of non-inferred gates: 0
  // ILP vars: 1675/1675
  // type: INFERRED
  // marked bad? no

  DFFQ_X1M_A12TR c0sm_b0m_v0m_tail_reg_0_ (.CK(clk), .Q(c0sm_b0m_v0m_tail_0_), .D(c0sm_b0m_v0m_n277));
  DFFQ_X1M_A12TR c0sm_b0m_v0m_tail_reg_1_ (.CK(clk), .Q(c0sm_b0m_v0m_tail_1_), .D(c0sm_b0m_v0m_n278));
endmodule
